
//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ../td_ccore_solutions/Connections__InBlocking_SysPE__InputType_Connections__SYN_--_134108c48ee88347694fbbe76a2ae1cc6142_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Sun May  3 14:21:41 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  mgc_out_dreg_v2 #(.rscid(32'sd1),
  .width(32'sd8)) data_rsci (
      .d(nl_data_rsci_d[7:0]),
      .z(data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd216),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__InBlocking_SysPE__AccumType_Connections__SYN_--_825475bfda2a8d92d42aecf1ac6780716115_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Sun May  3 14:21:38 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [31:0] this_msg;
  output [31:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  mgc_out_dreg_v2 #(.rscid(32'sd4),
  .width(32'sd32)) data_rsci (
      .d(nl_data_rsci_d[31:0]),
      .z(data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd215),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [31:0] this_msg;
  output [31:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ../td_ccore_solutions/Connections__OutBlocking_SysPE__InputType_Connections__SYN--_402b1caf9f8ccdd7cb3d4b7d690caecb5c96_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Sun May  3 14:21:35 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [7:0] this_msg;
  reg [7:0] this_msg;
  input [7:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [7:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd7),
  .width(32'sd8)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd214),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd218)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 8'b00000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_msg <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [7:0] this_msg;
  input [7:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__OutBlocking_SysPE__AccumType_Connections__SYN--_e8bd1f99c97a28ffba001f7e6172d9185bea_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Sun May  3 14:21:31 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [31:0] this_msg;
  reg [31:0] this_msg;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [31:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd8),
  .width(32'sd32)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd213),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd217)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_msg <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [31:0] this_msg;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_SysPE__InputType_Connections__S--_3a7d47f76e133e87373796c2bf8aa2f0618f_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Sun May  3 14:21:28 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB_core
    (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  mgc_out_dreg_v2 #(.rscid(32'sd15),
  .width(32'sd8)) data_rsci (
      .d(nl_data_rsci_d[7:0]),
      .z(data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd16),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd212),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB_core Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_SysPE__AccumType_Connections__S--_cf9160d9abd7b1b11f697cebc35a1c465d23_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Sun May  3 14:21:25 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB_core
// ------------------------------------------------------------------


module Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB_core
    (
  this_val, this_rdy, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  mgc_out_dreg_v2 #(.rscid(32'sd18),
  .width(32'sd1)) return_rsci (
      .d(this_rdy),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd211),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_val <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB
// ------------------------------------------------------------------


module Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk,
      ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [31:0] this_msg;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB_core Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
  assign this_msg = 32'b00000000000000000000000000000000;
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Sun May  3 14:22:03 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SysArray_AccumInRun_AccumInRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysArray_AccumInRun_AccumInRun_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysArray_AccumInRun_AccumInRun_fsm_1
  parameter
    AccumInRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysArray_AccumInRun_AccumInRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // AccumInRun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= AccumInRun_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_ActOutRun_ActOutRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysArray_ActOutRun_ActOutRun_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysArray_ActOutRun_ActOutRun_fsm_1
  parameter
    ActOutRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysArray_ActOutRun_ActOutRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // ActOutRun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= ActOutRun_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_WeightOutRun_WeightOutRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysArray_WeightOutRun_WeightOutRun_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysArray_WeightOutRun_WeightOutRun_fsm_1
  parameter
    WeightOutRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysArray_WeightOutRun_WeightOutRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // WeightOutRun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= WeightOutRun_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_PERun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysPE_PERun_PERun_fsm (
  clk, rst, PERun_wen, fsm_output
);
  input clk;
  input rst;
  input PERun_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysPE_PERun_PERun_fsm_1
  parameter
    PERun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysPE_PERun_PERun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // PERun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PERun_rlp_C_0;
    end
    else if ( PERun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_staller
// ------------------------------------------------------------------


module SysPE_PERun_staller (
  clk, rst, PERun_wen, PERun_wten, act_out_Push_mioi_wen_comp, accum_out_Push_mioi_wen_comp,
      weight_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PERun_wen;
  output PERun_wten;
  input act_out_Push_mioi_wen_comp;
  input accum_out_Push_mioi_wen_comp;
  input weight_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PERun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PERun_wen = act_out_Push_mioi_wen_comp & accum_out_Push_mioi_wen_comp &
      weight_out_Push_mioi_wen_comp;
  assign PERun_wten = PERun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PERun_wten_reg <= 1'b0;
    end
    else begin
      PERun_wten_reg <= ~ PERun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_out_Push_mioi_weight_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_weight_out_Push_mioi_weight_out_Push_mio_wait_dp (
  clk, rst, weight_out_Push_mioi_oswt, weight_out_Push_mioi_wen_comp, weight_out_Push_mioi_biwt,
      weight_out_Push_mioi_bdwt, weight_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input weight_out_Push_mioi_oswt;
  output weight_out_Push_mioi_wen_comp;
  input weight_out_Push_mioi_biwt;
  input weight_out_Push_mioi_bdwt;
  output weight_out_Push_mioi_bcwt;
  reg weight_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign weight_out_Push_mioi_wen_comp = (~ weight_out_Push_mioi_oswt) | weight_out_Push_mioi_biwt
      | weight_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      weight_out_Push_mioi_bcwt <= ~((~(weight_out_Push_mioi_bcwt | weight_out_Push_mioi_biwt))
          | weight_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_out_Push_mioi_weight_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_weight_out_Push_mioi_weight_out_Push_mio_wait_ctrl (
  PERun_wen, weight_out_Push_mioi_oswt, weight_out_Push_mioi_biwt, weight_out_Push_mioi_bdwt,
      weight_out_Push_mioi_bcwt, weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct,
      weight_out_Push_mioi_ccs_ccore_done_sync_vld, weight_out_Push_mioi_oswt_pff
);
  input PERun_wen;
  input weight_out_Push_mioi_oswt;
  output weight_out_Push_mioi_biwt;
  output weight_out_Push_mioi_bdwt;
  input weight_out_Push_mioi_bcwt;
  output weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input weight_out_Push_mioi_ccs_ccore_done_sync_vld;
  input weight_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign weight_out_Push_mioi_bdwt = weight_out_Push_mioi_oswt & PERun_wen;
  assign weight_out_Push_mioi_biwt = weight_out_Push_mioi_oswt & (~ weight_out_Push_mioi_bcwt)
      & weight_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct = weight_out_Push_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp (
  clk, rst, accum_out_Push_mioi_oswt, accum_out_Push_mioi_wen_comp, accum_out_Push_mioi_biwt,
      accum_out_Push_mioi_bdwt, accum_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_wen_comp;
  input accum_out_Push_mioi_biwt;
  input accum_out_Push_mioi_bdwt;
  output accum_out_Push_mioi_bcwt;
  reg accum_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign accum_out_Push_mioi_wen_comp = (~ accum_out_Push_mioi_oswt) | accum_out_Push_mioi_biwt
      | accum_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      accum_out_Push_mioi_bcwt <= ~((~(accum_out_Push_mioi_bcwt | accum_out_Push_mioi_biwt))
          | accum_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl (
  PERun_wen, accum_out_Push_mioi_oswt, accum_out_Push_mioi_biwt, accum_out_Push_mioi_bdwt,
      accum_out_Push_mioi_bcwt, accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct,
      accum_out_Push_mioi_ccs_ccore_done_sync_vld, accum_out_Push_mioi_oswt_pff
);
  input PERun_wen;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_biwt;
  output accum_out_Push_mioi_bdwt;
  input accum_out_Push_mioi_bcwt;
  output accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input accum_out_Push_mioi_ccs_ccore_done_sync_vld;
  input accum_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accum_out_Push_mioi_bdwt = accum_out_Push_mioi_oswt & PERun_wen;
  assign accum_out_Push_mioi_biwt = accum_out_Push_mioi_oswt & (~ accum_out_Push_mioi_bcwt)
      & accum_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct = accum_out_Push_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp (
  clk, rst, act_out_Push_mioi_oswt, act_out_Push_mioi_wen_comp, act_out_Push_mioi_biwt,
      act_out_Push_mioi_bdwt, act_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_wen_comp;
  input act_out_Push_mioi_biwt;
  input act_out_Push_mioi_bdwt;
  output act_out_Push_mioi_bcwt;
  reg act_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_out_Push_mioi_wen_comp = (~ act_out_Push_mioi_oswt) | act_out_Push_mioi_biwt
      | act_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_out_Push_mioi_bcwt <= ~((~(act_out_Push_mioi_bcwt | act_out_Push_mioi_biwt))
          | act_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl (
  PERun_wen, act_out_Push_mioi_oswt, act_out_Push_mioi_biwt, act_out_Push_mioi_bdwt,
      act_out_Push_mioi_bcwt, act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct,
      act_out_Push_mioi_ccs_ccore_done_sync_vld, act_out_Push_mioi_oswt_pff
);
  input PERun_wen;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_biwt;
  output act_out_Push_mioi_bdwt;
  input act_out_Push_mioi_bcwt;
  output act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input act_out_Push_mioi_ccs_ccore_done_sync_vld;
  input act_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_out_Push_mioi_bdwt = act_out_Push_mioi_oswt & PERun_wen;
  assign act_out_Push_mioi_biwt = act_out_Push_mioi_oswt & (~ act_out_Push_mioi_bcwt)
      & act_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct = act_out_Push_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp (
  clk, rst, accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_in_PopNB_mioi_return_rsc_z_mxwt,
      accum_in_PopNB_mioi_data_rsc_z, accum_in_PopNB_mioi_biwt, accum_in_PopNB_mioi_bdwt,
      accum_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  output accum_in_PopNB_mioi_return_rsc_z_mxwt;
  input [31:0] accum_in_PopNB_mioi_data_rsc_z;
  input accum_in_PopNB_mioi_biwt;
  input accum_in_PopNB_mioi_bdwt;
  input accum_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg accum_in_PopNB_mioi_bcwt;
  reg [31:0] accum_in_PopNB_mioi_data_rsc_z_bfwt;
  reg accum_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accum_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_32_2_2(accum_in_PopNB_mioi_data_rsc_z,
      accum_in_PopNB_mioi_data_rsc_z_bfwt, accum_in_PopNB_mioi_bcwt);
  assign accum_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(accum_in_PopNB_mioi_return_rsc_z,
      accum_in_PopNB_mioi_return_rsc_z_bfwt, accum_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_in_PopNB_mioi_bcwt <= 1'b0;
      accum_in_PopNB_mioi_data_rsc_z_bfwt <= 32'b00000000000000000000000000000000;
      accum_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      accum_in_PopNB_mioi_bcwt <= ~((~(accum_in_PopNB_mioi_bcwt | accum_in_PopNB_mioi_biwt))
          | accum_in_PopNB_mioi_bdwt);
      accum_in_PopNB_mioi_data_rsc_z_bfwt <= accum_in_PopNB_mioi_data_rsc_z_mxwt;
      accum_in_PopNB_mioi_return_rsc_z_bfwt <= accum_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl (
  PERun_wen, PERun_wten, accum_in_PopNB_mioi_oswt, accum_in_PopNB_mioi_biwt, accum_in_PopNB_mioi_bdwt,
      accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct, accum_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input PERun_wten;
  input accum_in_PopNB_mioi_oswt;
  output accum_in_PopNB_mioi_biwt;
  output accum_in_PopNB_mioi_bdwt;
  output accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input accum_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accum_in_PopNB_mioi_bdwt = accum_in_PopNB_mioi_oswt & PERun_wen;
  assign accum_in_PopNB_mioi_biwt = (~ PERun_wten) & accum_in_PopNB_mioi_oswt;
  assign accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct = accum_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp (
  clk, rst, act_in_PopNB_mioi_data_rsc_z_mxwt, act_in_PopNB_mioi_return_rsc_z_mxwt,
      act_in_PopNB_mioi_data_rsc_z, act_in_PopNB_mioi_biwt, act_in_PopNB_mioi_bdwt,
      act_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  output act_in_PopNB_mioi_return_rsc_z_mxwt;
  input [7:0] act_in_PopNB_mioi_data_rsc_z;
  input act_in_PopNB_mioi_biwt;
  input act_in_PopNB_mioi_bdwt;
  input act_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg act_in_PopNB_mioi_bcwt;
  reg [7:0] act_in_PopNB_mioi_data_rsc_z_bfwt;
  reg act_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign act_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_8_2_2(act_in_PopNB_mioi_data_rsc_z,
      act_in_PopNB_mioi_data_rsc_z_bfwt, act_in_PopNB_mioi_bcwt);
  assign act_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(act_in_PopNB_mioi_return_rsc_z,
      act_in_PopNB_mioi_return_rsc_z_bfwt, act_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_PopNB_mioi_bcwt <= 1'b0;
      act_in_PopNB_mioi_data_rsc_z_bfwt <= 8'b00000000;
      act_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      act_in_PopNB_mioi_bcwt <= ~((~(act_in_PopNB_mioi_bcwt | act_in_PopNB_mioi_biwt))
          | act_in_PopNB_mioi_bdwt);
      act_in_PopNB_mioi_data_rsc_z_bfwt <= act_in_PopNB_mioi_data_rsc_z_mxwt;
      act_in_PopNB_mioi_return_rsc_z_bfwt <= act_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl (
  PERun_wen, PERun_wten, act_in_PopNB_mioi_oswt, act_in_PopNB_mioi_biwt, act_in_PopNB_mioi_bdwt,
      act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct, act_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input PERun_wten;
  input act_in_PopNB_mioi_oswt;
  output act_in_PopNB_mioi_biwt;
  output act_in_PopNB_mioi_bdwt;
  output act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input act_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_PopNB_mioi_bdwt = act_in_PopNB_mioi_oswt & PERun_wen;
  assign act_in_PopNB_mioi_biwt = (~ PERun_wten) & act_in_PopNB_mioi_oswt;
  assign act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct = act_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp (
  clk, rst, weight_in_PopNB_mioi_data_rsc_z_mxwt, weight_in_PopNB_mioi_return_rsc_z_mxwt,
      weight_in_PopNB_mioi_data_rsc_z, weight_in_PopNB_mioi_biwt, weight_in_PopNB_mioi_bdwt,
      weight_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  output weight_in_PopNB_mioi_return_rsc_z_mxwt;
  input [7:0] weight_in_PopNB_mioi_data_rsc_z;
  input weight_in_PopNB_mioi_biwt;
  input weight_in_PopNB_mioi_bdwt;
  input weight_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg weight_in_PopNB_mioi_bcwt;
  reg [7:0] weight_in_PopNB_mioi_data_rsc_z_bfwt;
  reg weight_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign weight_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_8_2_2(weight_in_PopNB_mioi_data_rsc_z,
      weight_in_PopNB_mioi_data_rsc_z_bfwt, weight_in_PopNB_mioi_bcwt);
  assign weight_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(weight_in_PopNB_mioi_return_rsc_z,
      weight_in_PopNB_mioi_return_rsc_z_bfwt, weight_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_in_PopNB_mioi_bcwt <= 1'b0;
      weight_in_PopNB_mioi_data_rsc_z_bfwt <= 8'b00000000;
      weight_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      weight_in_PopNB_mioi_bcwt <= ~((~(weight_in_PopNB_mioi_bcwt | weight_in_PopNB_mioi_biwt))
          | weight_in_PopNB_mioi_bdwt);
      weight_in_PopNB_mioi_data_rsc_z_bfwt <= weight_in_PopNB_mioi_data_rsc_z_mxwt;
      weight_in_PopNB_mioi_return_rsc_z_bfwt <= weight_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl (
  PERun_wen, weight_in_PopNB_mioi_oswt, PERun_wten, weight_in_PopNB_mioi_biwt, weight_in_PopNB_mioi_bdwt,
      weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct, weight_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input weight_in_PopNB_mioi_oswt;
  input PERun_wten;
  output weight_in_PopNB_mioi_biwt;
  output weight_in_PopNB_mioi_bdwt;
  output weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input weight_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign weight_in_PopNB_mioi_bdwt = weight_in_PopNB_mioi_oswt & PERun_wen;
  assign weight_in_PopNB_mioi_biwt = (~ PERun_wten) & weight_in_PopNB_mioi_oswt;
  assign weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct = weight_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_AccumInRun
// ------------------------------------------------------------------


module SysArray_AccumInRun (
  clk, rst, accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_pff
);
  input clk;
  input rst;
  output accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_pff;


  // Interconnect Declarations
  wire [1:0] fsm_output;

  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_1;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_2;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_3;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_4;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_5;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_6;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_7;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7;

  // Interconnect Declarations for Component Instantiations 
  SysArray_AccumInRun_AccumInRun_fsm SysArray_AccumInRun_AccumInRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign p0_Unreachable_virtual_function_in_abstract_class_prb = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb  -> p0_Unreachable_virtual_function_in_abstract_class_prb );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_1 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_1 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1  -> p0_Unreachable_virtual_function_in_abstract_class_prb_1 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_2 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_2 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2  -> p0_Unreachable_virtual_function_in_abstract_class_prb_2 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_3 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_3 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3  -> p0_Unreachable_virtual_function_in_abstract_class_prb_3 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_4 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_4 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4  -> p0_Unreachable_virtual_function_in_abstract_class_prb_4 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_5 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_5 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5  -> p0_Unreachable_virtual_function_in_abstract_class_prb_5 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_6 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_6 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6  -> p0_Unreachable_virtual_function_in_abstract_class_prb_6 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_7 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_7 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7  -> p0_Unreachable_virtual_function_in_abstract_class_prb_7 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7 = 1'b0;
  assign accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_pff = fsm_output[1];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_ActOutRun
// ------------------------------------------------------------------


module SysArray_ActOutRun (
  clk, rst, act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_pff
);
  input clk;
  input rst;
  output act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_pff;


  // Interconnect Declarations
  wire [1:0] fsm_output;


  // Interconnect Declarations for Component Instantiations 
  SysArray_ActOutRun_ActOutRun_fsm SysArray_ActOutRun_ActOutRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_pff = fsm_output[1];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_WeightOutRun
// ------------------------------------------------------------------


module SysArray_WeightOutRun (
  clk, rst, weight_inter_7_0_val, weight_inter_7_1_val, weight_inter_7_2_val, weight_inter_7_3_val,
      weight_inter_7_4_val, weight_inter_7_5_val, weight_inter_7_6_val, weight_inter_7_7_val,
      weight_inter_7_0_rdy, weight_inter_7_1_rdy, weight_inter_7_2_rdy, weight_inter_7_3_rdy,
      weight_inter_7_4_rdy, weight_inter_7_5_rdy, weight_inter_7_6_rdy, weight_inter_7_7_rdy,
      weight_inter_7_0_msg, weight_inter_7_1_msg, weight_inter_7_2_msg, weight_inter_7_3_msg,
      weight_inter_7_4_msg, weight_inter_7_5_msg, weight_inter_7_6_msg, weight_inter_7_7_msg
);
  input clk;
  input rst;
  input weight_inter_7_0_val;
  input weight_inter_7_1_val;
  input weight_inter_7_2_val;
  input weight_inter_7_3_val;
  input weight_inter_7_4_val;
  input weight_inter_7_5_val;
  input weight_inter_7_6_val;
  input weight_inter_7_7_val;
  output weight_inter_7_0_rdy;
  output weight_inter_7_1_rdy;
  output weight_inter_7_2_rdy;
  output weight_inter_7_3_rdy;
  output weight_inter_7_4_rdy;
  output weight_inter_7_5_rdy;
  output weight_inter_7_6_rdy;
  output weight_inter_7_7_rdy;
  input [7:0] weight_inter_7_0_msg;
  input [7:0] weight_inter_7_1_msg;
  input [7:0] weight_inter_7_2_msg;
  input [7:0] weight_inter_7_3_msg;
  input [7:0] weight_inter_7_4_msg;
  input [7:0] weight_inter_7_5_msg;
  input [7:0] weight_inter_7_6_msg;
  input [7:0] weight_inter_7_7_msg;


  // Interconnect Declarations
  wire [7:0] weight_inter_PopNB_56_mioi_data_rsc_z;
  wire weight_inter_PopNB_56_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_57_mioi_data_rsc_z;
  wire weight_inter_PopNB_57_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_58_mioi_data_rsc_z;
  wire weight_inter_PopNB_58_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_59_mioi_data_rsc_z;
  wire weight_inter_PopNB_59_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_60_mioi_data_rsc_z;
  wire weight_inter_PopNB_60_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_61_mioi_data_rsc_z;
  wire weight_inter_PopNB_61_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_62_mioi_data_rsc_z;
  wire weight_inter_PopNB_62_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_63_mioi_data_rsc_z;
  wire weight_inter_PopNB_63_mioi_return_rsc_z;
  wire [1:0] fsm_output;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat;
  assign nl_weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat = fsm_output[1];
  wire [0:0] nl_weight_inter_PopNB_57_mioi_ccs_ccore_start_rsc_dat;
  assign nl_weight_inter_PopNB_57_mioi_ccs_ccore_start_rsc_dat = fsm_output[1];
  wire [0:0] nl_weight_inter_PopNB_58_mioi_ccs_ccore_start_rsc_dat;
  assign nl_weight_inter_PopNB_58_mioi_ccs_ccore_start_rsc_dat = fsm_output[1];
  wire [0:0] nl_weight_inter_PopNB_59_mioi_ccs_ccore_start_rsc_dat;
  assign nl_weight_inter_PopNB_59_mioi_ccs_ccore_start_rsc_dat = fsm_output[1];
  wire [0:0] nl_weight_inter_PopNB_60_mioi_ccs_ccore_start_rsc_dat;
  assign nl_weight_inter_PopNB_60_mioi_ccs_ccore_start_rsc_dat = fsm_output[1];
  wire [0:0] nl_weight_inter_PopNB_61_mioi_ccs_ccore_start_rsc_dat;
  assign nl_weight_inter_PopNB_61_mioi_ccs_ccore_start_rsc_dat = fsm_output[1];
  wire [0:0] nl_weight_inter_PopNB_62_mioi_ccs_ccore_start_rsc_dat;
  assign nl_weight_inter_PopNB_62_mioi_ccs_ccore_start_rsc_dat = fsm_output[1];
  wire [0:0] nl_weight_inter_PopNB_63_mioi_ccs_ccore_start_rsc_dat;
  assign nl_weight_inter_PopNB_63_mioi_ccs_ccore_start_rsc_dat = fsm_output[1];
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_56_mioi
      (
      .this_val(weight_inter_7_0_val),
      .this_rdy(weight_inter_7_0_rdy),
      .this_msg(weight_inter_7_0_msg),
      .data_rsc_z(weight_inter_PopNB_56_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_56_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(nl_weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat[0:0])
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_57_mioi
      (
      .this_val(weight_inter_7_1_val),
      .this_rdy(weight_inter_7_1_rdy),
      .this_msg(weight_inter_7_1_msg),
      .data_rsc_z(weight_inter_PopNB_57_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_57_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(nl_weight_inter_PopNB_57_mioi_ccs_ccore_start_rsc_dat[0:0])
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_58_mioi
      (
      .this_val(weight_inter_7_2_val),
      .this_rdy(weight_inter_7_2_rdy),
      .this_msg(weight_inter_7_2_msg),
      .data_rsc_z(weight_inter_PopNB_58_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_58_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(nl_weight_inter_PopNB_58_mioi_ccs_ccore_start_rsc_dat[0:0])
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_59_mioi
      (
      .this_val(weight_inter_7_3_val),
      .this_rdy(weight_inter_7_3_rdy),
      .this_msg(weight_inter_7_3_msg),
      .data_rsc_z(weight_inter_PopNB_59_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_59_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(nl_weight_inter_PopNB_59_mioi_ccs_ccore_start_rsc_dat[0:0])
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_60_mioi
      (
      .this_val(weight_inter_7_4_val),
      .this_rdy(weight_inter_7_4_rdy),
      .this_msg(weight_inter_7_4_msg),
      .data_rsc_z(weight_inter_PopNB_60_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_60_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(nl_weight_inter_PopNB_60_mioi_ccs_ccore_start_rsc_dat[0:0])
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_61_mioi
      (
      .this_val(weight_inter_7_5_val),
      .this_rdy(weight_inter_7_5_rdy),
      .this_msg(weight_inter_7_5_msg),
      .data_rsc_z(weight_inter_PopNB_61_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_61_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(nl_weight_inter_PopNB_61_mioi_ccs_ccore_start_rsc_dat[0:0])
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_62_mioi
      (
      .this_val(weight_inter_7_6_val),
      .this_rdy(weight_inter_7_6_rdy),
      .this_msg(weight_inter_7_6_msg),
      .data_rsc_z(weight_inter_PopNB_62_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_62_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(nl_weight_inter_PopNB_62_mioi_ccs_ccore_start_rsc_dat[0:0])
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_63_mioi
      (
      .this_val(weight_inter_7_7_val),
      .this_rdy(weight_inter_7_7_rdy),
      .this_msg(weight_inter_7_7_msg),
      .data_rsc_z(weight_inter_PopNB_63_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_63_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(nl_weight_inter_PopNB_63_mioi_ccs_ccore_start_rsc_dat[0:0])
    );
  SysArray_WeightOutRun_WeightOutRun_fsm SysArray_WeightOutRun_WeightOutRun_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_out_Push_mioi
// ------------------------------------------------------------------


module SysPE_PERun_weight_out_Push_mioi (
  clk, rst, weight_out_val, weight_out_rdy, weight_out_msg, PERun_wen, weight_out_Push_mioi_oswt,
      weight_out_Push_mioi_wen_comp, weight_out_Push_mioi_m_rsc_dat_PERun, weight_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;
  input PERun_wen;
  input weight_out_Push_mioi_oswt;
  output weight_out_Push_mioi_wen_comp;
  input [7:0] weight_out_Push_mioi_m_rsc_dat_PERun;
  input weight_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire weight_out_Push_mioi_biwt;
  wire weight_out_Push_mioi_bdwt;
  wire weight_out_Push_mioi_bcwt;
  wire weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  wire weight_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  weight_out_Push_mioi
      (
      .this_val(weight_out_val),
      .this_rdy(weight_out_rdy),
      .this_msg(weight_out_msg),
      .m_rsc_dat(weight_out_Push_mioi_m_rsc_dat_PERun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .ccs_ccore_done_sync_vld(weight_out_Push_mioi_ccs_ccore_done_sync_vld)
    );
  SysPE_PERun_weight_out_Push_mioi_weight_out_Push_mio_wait_ctrl SysPE_PERun_weight_out_Push_mioi_weight_out_Push_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .weight_out_Push_mioi_oswt(weight_out_Push_mioi_oswt),
      .weight_out_Push_mioi_biwt(weight_out_Push_mioi_biwt),
      .weight_out_Push_mioi_bdwt(weight_out_Push_mioi_bdwt),
      .weight_out_Push_mioi_bcwt(weight_out_Push_mioi_bcwt),
      .weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct(weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .weight_out_Push_mioi_ccs_ccore_done_sync_vld(weight_out_Push_mioi_ccs_ccore_done_sync_vld),
      .weight_out_Push_mioi_oswt_pff(weight_out_Push_mioi_oswt_pff)
    );
  SysPE_PERun_weight_out_Push_mioi_weight_out_Push_mio_wait_dp SysPE_PERun_weight_out_Push_mioi_weight_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .weight_out_Push_mioi_oswt(weight_out_Push_mioi_oswt),
      .weight_out_Push_mioi_wen_comp(weight_out_Push_mioi_wen_comp),
      .weight_out_Push_mioi_biwt(weight_out_Push_mioi_biwt),
      .weight_out_Push_mioi_bdwt(weight_out_Push_mioi_bdwt),
      .weight_out_Push_mioi_bcwt(weight_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi (
  clk, rst, accum_out_val, accum_out_rdy, accum_out_msg, PERun_wen, accum_out_Push_mioi_oswt,
      accum_out_Push_mioi_wen_comp, accum_out_Push_mioi_m_rsc_dat_PERun, accum_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;
  input PERun_wen;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_wen_comp;
  input [31:0] accum_out_Push_mioi_m_rsc_dat_PERun;
  input accum_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire accum_out_Push_mioi_biwt;
  wire accum_out_Push_mioi_bdwt;
  wire accum_out_Push_mioi_bcwt;
  wire accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  wire accum_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push  accum_out_Push_mioi
      (
      .this_val(accum_out_val),
      .this_rdy(accum_out_rdy),
      .this_msg(accum_out_msg),
      .m_rsc_dat(accum_out_Push_mioi_m_rsc_dat_PERun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .ccs_ccore_done_sync_vld(accum_out_Push_mioi_ccs_ccore_done_sync_vld)
    );
  SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .accum_out_Push_mioi_oswt(accum_out_Push_mioi_oswt),
      .accum_out_Push_mioi_biwt(accum_out_Push_mioi_biwt),
      .accum_out_Push_mioi_bdwt(accum_out_Push_mioi_bdwt),
      .accum_out_Push_mioi_bcwt(accum_out_Push_mioi_bcwt),
      .accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct(accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .accum_out_Push_mioi_ccs_ccore_done_sync_vld(accum_out_Push_mioi_ccs_ccore_done_sync_vld),
      .accum_out_Push_mioi_oswt_pff(accum_out_Push_mioi_oswt_pff)
    );
  SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .accum_out_Push_mioi_oswt(accum_out_Push_mioi_oswt),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_biwt(accum_out_Push_mioi_biwt),
      .accum_out_Push_mioi_bdwt(accum_out_Push_mioi_bdwt),
      .accum_out_Push_mioi_bcwt(accum_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi (
  clk, rst, act_out_val, act_out_rdy, act_out_msg, PERun_wen, act_out_Push_mioi_oswt,
      act_out_Push_mioi_wen_comp, act_out_Push_mioi_m_rsc_dat_PERun, act_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  input PERun_wen;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_wen_comp;
  input [7:0] act_out_Push_mioi_m_rsc_dat_PERun;
  input act_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_out_Push_mioi_biwt;
  wire act_out_Push_mioi_bdwt;
  wire act_out_Push_mioi_bcwt;
  wire act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  wire act_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_out_Push_mioi
      (
      .this_val(act_out_val),
      .this_rdy(act_out_rdy),
      .this_msg(act_out_msg),
      .m_rsc_dat(act_out_Push_mioi_m_rsc_dat_PERun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .ccs_ccore_done_sync_vld(act_out_Push_mioi_ccs_ccore_done_sync_vld)
    );
  SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .act_out_Push_mioi_oswt(act_out_Push_mioi_oswt),
      .act_out_Push_mioi_biwt(act_out_Push_mioi_biwt),
      .act_out_Push_mioi_bdwt(act_out_Push_mioi_bdwt),
      .act_out_Push_mioi_bcwt(act_out_Push_mioi_bcwt),
      .act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct(act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .act_out_Push_mioi_ccs_ccore_done_sync_vld(act_out_Push_mioi_ccs_ccore_done_sync_vld),
      .act_out_Push_mioi_oswt_pff(act_out_Push_mioi_oswt_pff)
    );
  SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_out_Push_mioi_oswt(act_out_Push_mioi_oswt),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .act_out_Push_mioi_biwt(act_out_Push_mioi_biwt),
      .act_out_Push_mioi_bdwt(act_out_Push_mioi_bdwt),
      .act_out_Push_mioi_bcwt(act_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi (
  clk, rst, accum_in_val, accum_in_rdy, accum_in_msg, PERun_wen, PERun_wten, accum_in_PopNB_mioi_oswt,
      accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_in_PopNB_mioi_return_rsc_z_mxwt,
      accum_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  input PERun_wen;
  input PERun_wten;
  input accum_in_PopNB_mioi_oswt;
  output [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  output accum_in_PopNB_mioi_return_rsc_z_mxwt;
  input accum_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [31:0] accum_in_PopNB_mioi_data_rsc_z;
  wire accum_in_PopNB_mioi_biwt;
  wire accum_in_PopNB_mioi_bdwt;
  wire accum_in_PopNB_mioi_return_rsc_z;
  wire accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB  accum_in_PopNB_mioi
      (
      .this_val(accum_in_val),
      .this_rdy(accum_in_rdy),
      .this_msg(accum_in_msg),
      .data_rsc_z(accum_in_PopNB_mioi_data_rsc_z),
      .return_rsc_z(accum_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
  SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .accum_in_PopNB_mioi_oswt(accum_in_PopNB_mioi_oswt),
      .accum_in_PopNB_mioi_biwt(accum_in_PopNB_mioi_biwt),
      .accum_in_PopNB_mioi_bdwt(accum_in_PopNB_mioi_bdwt),
      .accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct(accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .accum_in_PopNB_mioi_oswt_pff(accum_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .accum_in_PopNB_mioi_data_rsc_z_mxwt(accum_in_PopNB_mioi_data_rsc_z_mxwt),
      .accum_in_PopNB_mioi_return_rsc_z_mxwt(accum_in_PopNB_mioi_return_rsc_z_mxwt),
      .accum_in_PopNB_mioi_data_rsc_z(accum_in_PopNB_mioi_data_rsc_z),
      .accum_in_PopNB_mioi_biwt(accum_in_PopNB_mioi_biwt),
      .accum_in_PopNB_mioi_bdwt(accum_in_PopNB_mioi_bdwt),
      .accum_in_PopNB_mioi_return_rsc_z(accum_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi (
  clk, rst, act_in_val, act_in_rdy, act_in_msg, PERun_wen, PERun_wten, act_in_PopNB_mioi_oswt,
      act_in_PopNB_mioi_data_rsc_z_mxwt, act_in_PopNB_mioi_return_rsc_z_mxwt, act_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input PERun_wen;
  input PERun_wten;
  input act_in_PopNB_mioi_oswt;
  output [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  output act_in_PopNB_mioi_return_rsc_z_mxwt;
  input act_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [7:0] act_in_PopNB_mioi_data_rsc_z;
  wire act_in_PopNB_mioi_biwt;
  wire act_in_PopNB_mioi_bdwt;
  wire act_in_PopNB_mioi_return_rsc_z;
  wire act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB  act_in_PopNB_mioi
      (
      .this_val(act_in_val),
      .this_rdy(act_in_rdy),
      .this_msg(act_in_msg),
      .data_rsc_z(act_in_PopNB_mioi_data_rsc_z),
      .return_rsc_z(act_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
  SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_in_PopNB_mioi_oswt(act_in_PopNB_mioi_oswt),
      .act_in_PopNB_mioi_biwt(act_in_PopNB_mioi_biwt),
      .act_in_PopNB_mioi_bdwt(act_in_PopNB_mioi_bdwt),
      .act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct(act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .act_in_PopNB_mioi_oswt_pff(act_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_PopNB_mioi_data_rsc_z_mxwt(act_in_PopNB_mioi_data_rsc_z_mxwt),
      .act_in_PopNB_mioi_return_rsc_z_mxwt(act_in_PopNB_mioi_return_rsc_z_mxwt),
      .act_in_PopNB_mioi_data_rsc_z(act_in_PopNB_mioi_data_rsc_z),
      .act_in_PopNB_mioi_biwt(act_in_PopNB_mioi_biwt),
      .act_in_PopNB_mioi_bdwt(act_in_PopNB_mioi_bdwt),
      .act_in_PopNB_mioi_return_rsc_z(act_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, PERun_wen, weight_in_PopNB_mioi_oswt,
      PERun_wten, weight_in_PopNB_mioi_data_rsc_z_mxwt, weight_in_PopNB_mioi_return_rsc_z_mxwt,
      weight_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input PERun_wen;
  input weight_in_PopNB_mioi_oswt;
  input PERun_wten;
  output [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  output weight_in_PopNB_mioi_return_rsc_z_mxwt;
  input weight_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [7:0] weight_in_PopNB_mioi_data_rsc_z;
  wire weight_in_PopNB_mioi_biwt;
  wire weight_in_PopNB_mioi_bdwt;
  wire weight_in_PopNB_mioi_return_rsc_z;
  wire weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_in_PopNB_mioi
      (
      .this_val(weight_in_val),
      .this_rdy(weight_in_rdy),
      .this_msg(weight_in_msg),
      .data_rsc_z(weight_in_PopNB_mioi_data_rsc_z),
      .return_rsc_z(weight_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
  SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .weight_in_PopNB_mioi_oswt(weight_in_PopNB_mioi_oswt),
      .PERun_wten(PERun_wten),
      .weight_in_PopNB_mioi_biwt(weight_in_PopNB_mioi_biwt),
      .weight_in_PopNB_mioi_bdwt(weight_in_PopNB_mioi_bdwt),
      .weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct(weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .weight_in_PopNB_mioi_oswt_pff(weight_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .weight_in_PopNB_mioi_data_rsc_z_mxwt(weight_in_PopNB_mioi_data_rsc_z_mxwt),
      .weight_in_PopNB_mioi_return_rsc_z_mxwt(weight_in_PopNB_mioi_return_rsc_z_mxwt),
      .weight_in_PopNB_mioi_data_rsc_z(weight_in_PopNB_mioi_data_rsc_z),
      .weight_in_PopNB_mioi_biwt(weight_in_PopNB_mioi_biwt),
      .weight_in_PopNB_mioi_bdwt(weight_in_PopNB_mioi_bdwt),
      .weight_in_PopNB_mioi_return_rsc_z(weight_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun
// ------------------------------------------------------------------


module SysPE_PERun (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, act_in_val, act_in_rdy,
      act_in_msg, accum_in_val, accum_in_rdy, accum_in_msg, weight_out_val, weight_out_rdy,
      weight_out_msg, act_out_val, act_out_rdy, act_out_msg, accum_out_val, accum_out_rdy,
      accum_out_msg
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;


  // Interconnect Declarations
  wire PERun_wen;
  wire PERun_wten;
  wire [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  wire weight_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  wire act_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  wire accum_in_PopNB_mioi_return_rsc_z_mxwt;
  wire act_out_Push_mioi_wen_comp;
  wire accum_out_Push_mioi_wen_comp;
  wire weight_out_Push_mioi_wen_comp;
  wire [1:0] fsm_output;
  wire while_while_or_tmp;
  wire and_dcpl;
  wire is_accum_in_sva_dfm_1;
  reg is_accum_in_sva;
  reg is_act_in_sva;
  wire while_land_lpi_1_dfm_1;
  reg reg_weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  wire is_accum_in_63_and_cse;
  wire and_4_cse;
  wire mux_7_cse;
  wire and_9_rmff;
  wire and_7_rmff;
  wire and_2_rmff;
  reg [7:0] act_reg_sva;
  wire [7:0] act_out_Push_mioi_m_rsc_dat_PERun_mx1;
  reg [7:0] weight_reg_sva;
  wire [31:0] accum_reg_sva_mx0;
  reg [31:0] accum_reg_sva;

  wire[0:0] or_3_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_11_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] or_18_nl;
  wire[0:0] nor_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff;
  assign nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff =
      fsm_output[1];
  wire[0:0] or_nl;
  wire [7:0] nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun;
  assign or_nl = is_act_in_sva | (fsm_output[0]);
  assign nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun
      = MUX_v_8_2_2(act_in_PopNB_mioi_data_rsc_z_mxwt, act_reg_sva, or_nl);
  wire[15:0] while_if_3_accum_out_reg_mul_nl;
  wire[7:0] while_if_mux_1_nl;
  wire [31:0] nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun;
  assign while_if_mux_1_nl = MUX_v_8_2_2(weight_reg_sva, weight_in_PopNB_mioi_data_rsc_z_mxwt,
      weight_in_PopNB_mioi_return_rsc_z_mxwt);
  assign while_if_3_accum_out_reg_mul_nl = conv_s2u_16_16($signed((act_out_Push_mioi_m_rsc_dat_PERun_mx1))
      * $signed((while_if_mux_1_nl)));
  assign nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun
      = conv_s2u_16_32(while_if_3_accum_out_reg_mul_nl) + accum_reg_sva_mx0;
  wire [7:0] nl_SysPE_PERun_weight_out_Push_mioi_inst_weight_out_Push_mioi_m_rsc_dat_PERun;
  assign nl_SysPE_PERun_weight_out_Push_mioi_inst_weight_out_Push_mioi_m_rsc_dat_PERun
      = weight_reg_sva;
  SysPE_PERun_weight_in_PopNB_mioi SysPE_PERun_weight_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_val),
      .weight_in_rdy(weight_in_rdy),
      .weight_in_msg(weight_in_msg),
      .PERun_wen(PERun_wen),
      .weight_in_PopNB_mioi_oswt(reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .PERun_wten(PERun_wten),
      .weight_in_PopNB_mioi_data_rsc_z_mxwt(weight_in_PopNB_mioi_data_rsc_z_mxwt),
      .weight_in_PopNB_mioi_return_rsc_z_mxwt(weight_in_PopNB_mioi_return_rsc_z_mxwt),
      .weight_in_PopNB_mioi_oswt_pff(nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff[0:0])
    );
  SysPE_PERun_act_in_PopNB_mioi SysPE_PERun_act_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .act_in_val(act_in_val),
      .act_in_rdy(act_in_rdy),
      .act_in_msg(act_in_msg),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_in_PopNB_mioi_oswt(reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .act_in_PopNB_mioi_data_rsc_z_mxwt(act_in_PopNB_mioi_data_rsc_z_mxwt),
      .act_in_PopNB_mioi_return_rsc_z_mxwt(act_in_PopNB_mioi_return_rsc_z_mxwt),
      .act_in_PopNB_mioi_oswt_pff(and_9_rmff)
    );
  SysPE_PERun_accum_in_PopNB_mioi SysPE_PERun_accum_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .accum_in_val(accum_in_val),
      .accum_in_rdy(accum_in_rdy),
      .accum_in_msg(accum_in_msg),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .accum_in_PopNB_mioi_oswt(reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .accum_in_PopNB_mioi_data_rsc_z_mxwt(accum_in_PopNB_mioi_data_rsc_z_mxwt),
      .accum_in_PopNB_mioi_return_rsc_z_mxwt(accum_in_PopNB_mioi_return_rsc_z_mxwt),
      .accum_in_PopNB_mioi_oswt_pff(and_7_rmff)
    );
  SysPE_PERun_act_out_Push_mioi SysPE_PERun_act_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .act_out_val(act_out_val),
      .act_out_rdy(act_out_rdy),
      .act_out_msg(act_out_msg),
      .PERun_wen(PERun_wen),
      .act_out_Push_mioi_oswt(reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .act_out_Push_mioi_m_rsc_dat_PERun(nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun[7:0]),
      .act_out_Push_mioi_oswt_pff(and_4_cse)
    );
  SysPE_PERun_accum_out_Push_mioi SysPE_PERun_accum_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .accum_out_val(accum_out_val),
      .accum_out_rdy(accum_out_rdy),
      .accum_out_msg(accum_out_msg),
      .PERun_wen(PERun_wen),
      .accum_out_Push_mioi_oswt(reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_m_rsc_dat_PERun(nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun[31:0]),
      .accum_out_Push_mioi_oswt_pff(and_4_cse)
    );
  SysPE_PERun_weight_out_Push_mioi SysPE_PERun_weight_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .weight_out_val(weight_out_val),
      .weight_out_rdy(weight_out_rdy),
      .weight_out_msg(weight_out_msg),
      .PERun_wen(PERun_wen),
      .weight_out_Push_mioi_oswt(reg_weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .weight_out_Push_mioi_wen_comp(weight_out_Push_mioi_wen_comp),
      .weight_out_Push_mioi_m_rsc_dat_PERun(nl_SysPE_PERun_weight_out_Push_mioi_inst_weight_out_Push_mioi_m_rsc_dat_PERun[7:0]),
      .weight_out_Push_mioi_oswt_pff(and_2_rmff)
    );
  SysPE_PERun_staller SysPE_PERun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp),
      .weight_out_Push_mioi_wen_comp(weight_out_Push_mioi_wen_comp)
    );
  SysPE_PERun_PERun_fsm SysPE_PERun_PERun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PERun_wen(PERun_wen),
      .fsm_output(fsm_output)
    );
  assign and_2_rmff = weight_in_PopNB_mioi_return_rsc_z_mxwt & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  assign and_4_cse = and_dcpl & is_accum_in_sva_dfm_1;
  assign or_3_nl = (~ accum_in_PopNB_mioi_return_rsc_z_mxwt) | is_act_in_sva | act_in_PopNB_mioi_return_rsc_z_mxwt
      | (~ reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse);
  assign mux_7_cse = MUX_s_1_2_2((or_3_nl), and_dcpl, is_accum_in_sva);
  assign and_7_rmff = mux_7_cse & (fsm_output[1]);
  assign mux_8_nl = MUX_s_1_2_2(is_act_in_sva, while_while_or_tmp, reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse);
  assign or_11_nl = reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse
      | (~ is_act_in_sva);
  assign mux_9_nl = MUX_s_1_2_2((~ (mux_8_nl)), (or_11_nl), is_accum_in_sva_dfm_1);
  assign and_9_rmff = (mux_9_nl) & (fsm_output[1]);
  assign is_accum_in_63_and_cse = PERun_wen & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  assign act_out_Push_mioi_m_rsc_dat_PERun_mx1 = MUX_v_8_2_2(act_in_PopNB_mioi_data_rsc_z_mxwt,
      act_reg_sva, is_act_in_sva);
  assign accum_reg_sva_mx0 = MUX_v_32_2_2(accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_reg_sva,
      is_accum_in_sva);
  assign is_accum_in_sva_dfm_1 = accum_in_PopNB_mioi_return_rsc_z_mxwt | is_accum_in_sva;
  assign while_land_lpi_1_dfm_1 = is_accum_in_sva_dfm_1 & while_while_or_tmp;
  assign while_while_or_tmp = act_in_PopNB_mioi_return_rsc_z_mxwt | is_act_in_sva;
  assign and_dcpl = while_while_or_tmp & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
    end
    else if ( PERun_wen ) begin
      reg_weight_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_2_rmff;
      reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_4_cse;
      reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_7_rmff;
      reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_9_rmff;
      reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= fsm_output[1];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      is_accum_in_sva <= 1'b0;
      is_act_in_sva <= 1'b0;
    end
    else if ( is_accum_in_63_and_cse ) begin
      is_accum_in_sva <= is_accum_in_sva_dfm_1 & (~ while_land_lpi_1_dfm_1);
      is_act_in_sva <= while_while_or_tmp & (~ while_land_lpi_1_dfm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_reg_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( PERun_wen & (~ mux_7_cse) ) begin
      accum_reg_sva <= accum_reg_sva_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_reg_sva <= 8'b00000000;
    end
    else if ( PERun_wen & (mux_6_nl) ) begin
      act_reg_sva <= act_out_Push_mioi_m_rsc_dat_PERun_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_reg_sva <= 8'b00000000;
    end
    else if ( PERun_wen & weight_in_PopNB_mioi_return_rsc_z_mxwt & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse
        ) begin
      weight_reg_sva <= weight_in_PopNB_mioi_data_rsc_z_mxwt;
    end
  end
  assign or_18_nl = is_act_in_sva | (act_in_PopNB_mioi_return_rsc_z_mxwt & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse);
  assign nor_nl = ~((~ is_act_in_sva) | reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse);
  assign mux_6_nl = MUX_s_1_2_2((or_18_nl), (nor_nl), is_accum_in_sva_dfm_1);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [15:0] conv_s2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_16 = vector;
  end
  endfunction


  function automatic [31:0] conv_s2u_16_32 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_32 = {{16{vector[15]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE
// ------------------------------------------------------------------


module SysPE (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, act_in_val, act_in_rdy,
      act_in_msg, accum_in_val, accum_in_rdy, accum_in_msg, weight_out_val, weight_out_rdy,
      weight_out_msg, act_out_val, act_out_rdy, act_out_msg, accum_out_val, accum_out_rdy,
      accum_out_msg
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;



  // Interconnect Declarations for Component Instantiations 
  SysPE_PERun SysPE_PERun_inst (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_val),
      .weight_in_rdy(weight_in_rdy),
      .weight_in_msg(weight_in_msg),
      .act_in_val(act_in_val),
      .act_in_rdy(act_in_rdy),
      .act_in_msg(act_in_msg),
      .accum_in_val(accum_in_val),
      .accum_in_rdy(accum_in_rdy),
      .accum_in_msg(accum_in_msg),
      .weight_out_val(weight_out_val),
      .weight_out_rdy(weight_out_rdy),
      .weight_out_msg(weight_out_msg),
      .act_out_val(act_out_val),
      .act_out_rdy(act_out_rdy),
      .act_out_msg(act_out_msg),
      .accum_out_val(accum_out_val),
      .accum_out_rdy(accum_out_rdy),
      .accum_out_msg(accum_out_msg)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_rtl
// ------------------------------------------------------------------


module SysArray_rtl (
  clk, rst, weight_in_vec_0_val, weight_in_vec_1_val, weight_in_vec_2_val, weight_in_vec_3_val,
      weight_in_vec_4_val, weight_in_vec_5_val, weight_in_vec_6_val, weight_in_vec_7_val,
      weight_in_vec_0_rdy, weight_in_vec_1_rdy, weight_in_vec_2_rdy, weight_in_vec_3_rdy,
      weight_in_vec_4_rdy, weight_in_vec_5_rdy, weight_in_vec_6_rdy, weight_in_vec_7_rdy,
      weight_in_vec_0_msg, weight_in_vec_1_msg, weight_in_vec_2_msg, weight_in_vec_3_msg,
      weight_in_vec_4_msg, weight_in_vec_5_msg, weight_in_vec_6_msg, weight_in_vec_7_msg,
      act_in_vec_0_val, act_in_vec_1_val, act_in_vec_2_val, act_in_vec_3_val, act_in_vec_4_val,
      act_in_vec_5_val, act_in_vec_6_val, act_in_vec_7_val, act_in_vec_0_rdy, act_in_vec_1_rdy,
      act_in_vec_2_rdy, act_in_vec_3_rdy, act_in_vec_4_rdy, act_in_vec_5_rdy, act_in_vec_6_rdy,
      act_in_vec_7_rdy, act_in_vec_0_msg, act_in_vec_1_msg, act_in_vec_2_msg, act_in_vec_3_msg,
      act_in_vec_4_msg, act_in_vec_5_msg, act_in_vec_6_msg, act_in_vec_7_msg, accum_out_vec_0_val,
      accum_out_vec_1_val, accum_out_vec_2_val, accum_out_vec_3_val, accum_out_vec_4_val,
      accum_out_vec_5_val, accum_out_vec_6_val, accum_out_vec_7_val, accum_out_vec_0_rdy,
      accum_out_vec_1_rdy, accum_out_vec_2_rdy, accum_out_vec_3_rdy, accum_out_vec_4_rdy,
      accum_out_vec_5_rdy, accum_out_vec_6_rdy, accum_out_vec_7_rdy, accum_out_vec_0_msg,
      accum_out_vec_1_msg, accum_out_vec_2_msg, accum_out_vec_3_msg, accum_out_vec_4_msg,
      accum_out_vec_5_msg, accum_out_vec_6_msg, accum_out_vec_7_msg
);
  input clk;
  input rst;
  input weight_in_vec_0_val;
  input weight_in_vec_1_val;
  input weight_in_vec_2_val;
  input weight_in_vec_3_val;
  input weight_in_vec_4_val;
  input weight_in_vec_5_val;
  input weight_in_vec_6_val;
  input weight_in_vec_7_val;
  output weight_in_vec_0_rdy;
  output weight_in_vec_1_rdy;
  output weight_in_vec_2_rdy;
  output weight_in_vec_3_rdy;
  output weight_in_vec_4_rdy;
  output weight_in_vec_5_rdy;
  output weight_in_vec_6_rdy;
  output weight_in_vec_7_rdy;
  input [7:0] weight_in_vec_0_msg;
  input [7:0] weight_in_vec_1_msg;
  input [7:0] weight_in_vec_2_msg;
  input [7:0] weight_in_vec_3_msg;
  input [7:0] weight_in_vec_4_msg;
  input [7:0] weight_in_vec_5_msg;
  input [7:0] weight_in_vec_6_msg;
  input [7:0] weight_in_vec_7_msg;
  input act_in_vec_0_val;
  input act_in_vec_1_val;
  input act_in_vec_2_val;
  input act_in_vec_3_val;
  input act_in_vec_4_val;
  input act_in_vec_5_val;
  input act_in_vec_6_val;
  input act_in_vec_7_val;
  output act_in_vec_0_rdy;
  output act_in_vec_1_rdy;
  output act_in_vec_2_rdy;
  output act_in_vec_3_rdy;
  output act_in_vec_4_rdy;
  output act_in_vec_5_rdy;
  output act_in_vec_6_rdy;
  output act_in_vec_7_rdy;
  input [7:0] act_in_vec_0_msg;
  input [7:0] act_in_vec_1_msg;
  input [7:0] act_in_vec_2_msg;
  input [7:0] act_in_vec_3_msg;
  input [7:0] act_in_vec_4_msg;
  input [7:0] act_in_vec_5_msg;
  input [7:0] act_in_vec_6_msg;
  input [7:0] act_in_vec_7_msg;
  output accum_out_vec_0_val;
  output accum_out_vec_1_val;
  output accum_out_vec_2_val;
  output accum_out_vec_3_val;
  output accum_out_vec_4_val;
  output accum_out_vec_5_val;
  output accum_out_vec_6_val;
  output accum_out_vec_7_val;
  input accum_out_vec_0_rdy;
  input accum_out_vec_1_rdy;
  input accum_out_vec_2_rdy;
  input accum_out_vec_3_rdy;
  input accum_out_vec_4_rdy;
  input accum_out_vec_5_rdy;
  input accum_out_vec_6_rdy;
  input accum_out_vec_7_rdy;
  output [31:0] accum_out_vec_0_msg;
  output [31:0] accum_out_vec_1_msg;
  output [31:0] accum_out_vec_2_msg;
  output [31:0] accum_out_vec_3_msg;
  output [31:0] accum_out_vec_4_msg;
  output [31:0] accum_out_vec_5_msg;
  output [31:0] accum_out_vec_6_msg;
  output [31:0] accum_out_vec_7_msg;


  // Interconnect Declarations
  wire weight_inter_0_0_val;
  wire weight_inter_0_1_val;
  wire weight_inter_0_2_val;
  wire weight_inter_0_3_val;
  wire weight_inter_0_4_val;
  wire weight_inter_0_5_val;
  wire weight_inter_0_6_val;
  wire weight_inter_0_7_val;
  wire weight_inter_1_0_val;
  wire weight_inter_1_1_val;
  wire weight_inter_1_2_val;
  wire weight_inter_1_3_val;
  wire weight_inter_1_4_val;
  wire weight_inter_1_5_val;
  wire weight_inter_1_6_val;
  wire weight_inter_1_7_val;
  wire weight_inter_2_0_val;
  wire weight_inter_2_1_val;
  wire weight_inter_2_2_val;
  wire weight_inter_2_3_val;
  wire weight_inter_2_4_val;
  wire weight_inter_2_5_val;
  wire weight_inter_2_6_val;
  wire weight_inter_2_7_val;
  wire weight_inter_3_0_val;
  wire weight_inter_3_1_val;
  wire weight_inter_3_2_val;
  wire weight_inter_3_3_val;
  wire weight_inter_3_4_val;
  wire weight_inter_3_5_val;
  wire weight_inter_3_6_val;
  wire weight_inter_3_7_val;
  wire weight_inter_4_0_val;
  wire weight_inter_4_1_val;
  wire weight_inter_4_2_val;
  wire weight_inter_4_3_val;
  wire weight_inter_4_4_val;
  wire weight_inter_4_5_val;
  wire weight_inter_4_6_val;
  wire weight_inter_4_7_val;
  wire weight_inter_5_0_val;
  wire weight_inter_5_1_val;
  wire weight_inter_5_2_val;
  wire weight_inter_5_3_val;
  wire weight_inter_5_4_val;
  wire weight_inter_5_5_val;
  wire weight_inter_5_6_val;
  wire weight_inter_5_7_val;
  wire weight_inter_6_0_val;
  wire weight_inter_6_1_val;
  wire weight_inter_6_2_val;
  wire weight_inter_6_3_val;
  wire weight_inter_6_4_val;
  wire weight_inter_6_5_val;
  wire weight_inter_6_6_val;
  wire weight_inter_6_7_val;
  wire weight_inter_7_0_val;
  wire weight_inter_7_1_val;
  wire weight_inter_7_2_val;
  wire weight_inter_7_3_val;
  wire weight_inter_7_4_val;
  wire weight_inter_7_5_val;
  wire weight_inter_7_6_val;
  wire weight_inter_7_7_val;
  wire weight_inter_0_0_rdy;
  wire weight_inter_0_1_rdy;
  wire weight_inter_0_2_rdy;
  wire weight_inter_0_3_rdy;
  wire weight_inter_0_4_rdy;
  wire weight_inter_0_5_rdy;
  wire weight_inter_0_6_rdy;
  wire weight_inter_0_7_rdy;
  wire weight_inter_1_0_rdy;
  wire weight_inter_1_1_rdy;
  wire weight_inter_1_2_rdy;
  wire weight_inter_1_3_rdy;
  wire weight_inter_1_4_rdy;
  wire weight_inter_1_5_rdy;
  wire weight_inter_1_6_rdy;
  wire weight_inter_1_7_rdy;
  wire weight_inter_2_0_rdy;
  wire weight_inter_2_1_rdy;
  wire weight_inter_2_2_rdy;
  wire weight_inter_2_3_rdy;
  wire weight_inter_2_4_rdy;
  wire weight_inter_2_5_rdy;
  wire weight_inter_2_6_rdy;
  wire weight_inter_2_7_rdy;
  wire weight_inter_3_0_rdy;
  wire weight_inter_3_1_rdy;
  wire weight_inter_3_2_rdy;
  wire weight_inter_3_3_rdy;
  wire weight_inter_3_4_rdy;
  wire weight_inter_3_5_rdy;
  wire weight_inter_3_6_rdy;
  wire weight_inter_3_7_rdy;
  wire weight_inter_4_0_rdy;
  wire weight_inter_4_1_rdy;
  wire weight_inter_4_2_rdy;
  wire weight_inter_4_3_rdy;
  wire weight_inter_4_4_rdy;
  wire weight_inter_4_5_rdy;
  wire weight_inter_4_6_rdy;
  wire weight_inter_4_7_rdy;
  wire weight_inter_5_0_rdy;
  wire weight_inter_5_1_rdy;
  wire weight_inter_5_2_rdy;
  wire weight_inter_5_3_rdy;
  wire weight_inter_5_4_rdy;
  wire weight_inter_5_5_rdy;
  wire weight_inter_5_6_rdy;
  wire weight_inter_5_7_rdy;
  wire weight_inter_6_0_rdy;
  wire weight_inter_6_1_rdy;
  wire weight_inter_6_2_rdy;
  wire weight_inter_6_3_rdy;
  wire weight_inter_6_4_rdy;
  wire weight_inter_6_5_rdy;
  wire weight_inter_6_6_rdy;
  wire weight_inter_6_7_rdy;
  wire weight_inter_7_0_rdy;
  wire weight_inter_7_1_rdy;
  wire weight_inter_7_2_rdy;
  wire weight_inter_7_3_rdy;
  wire weight_inter_7_4_rdy;
  wire weight_inter_7_5_rdy;
  wire weight_inter_7_6_rdy;
  wire weight_inter_7_7_rdy;
  wire [7:0] weight_inter_0_0_msg;
  wire [7:0] weight_inter_0_1_msg;
  wire [7:0] weight_inter_0_2_msg;
  wire [7:0] weight_inter_0_3_msg;
  wire [7:0] weight_inter_0_4_msg;
  wire [7:0] weight_inter_0_5_msg;
  wire [7:0] weight_inter_0_6_msg;
  wire [7:0] weight_inter_0_7_msg;
  wire [7:0] weight_inter_1_0_msg;
  wire [7:0] weight_inter_1_1_msg;
  wire [7:0] weight_inter_1_2_msg;
  wire [7:0] weight_inter_1_3_msg;
  wire [7:0] weight_inter_1_4_msg;
  wire [7:0] weight_inter_1_5_msg;
  wire [7:0] weight_inter_1_6_msg;
  wire [7:0] weight_inter_1_7_msg;
  wire [7:0] weight_inter_2_0_msg;
  wire [7:0] weight_inter_2_1_msg;
  wire [7:0] weight_inter_2_2_msg;
  wire [7:0] weight_inter_2_3_msg;
  wire [7:0] weight_inter_2_4_msg;
  wire [7:0] weight_inter_2_5_msg;
  wire [7:0] weight_inter_2_6_msg;
  wire [7:0] weight_inter_2_7_msg;
  wire [7:0] weight_inter_3_0_msg;
  wire [7:0] weight_inter_3_1_msg;
  wire [7:0] weight_inter_3_2_msg;
  wire [7:0] weight_inter_3_3_msg;
  wire [7:0] weight_inter_3_4_msg;
  wire [7:0] weight_inter_3_5_msg;
  wire [7:0] weight_inter_3_6_msg;
  wire [7:0] weight_inter_3_7_msg;
  wire [7:0] weight_inter_4_0_msg;
  wire [7:0] weight_inter_4_1_msg;
  wire [7:0] weight_inter_4_2_msg;
  wire [7:0] weight_inter_4_3_msg;
  wire [7:0] weight_inter_4_4_msg;
  wire [7:0] weight_inter_4_5_msg;
  wire [7:0] weight_inter_4_6_msg;
  wire [7:0] weight_inter_4_7_msg;
  wire [7:0] weight_inter_5_0_msg;
  wire [7:0] weight_inter_5_1_msg;
  wire [7:0] weight_inter_5_2_msg;
  wire [7:0] weight_inter_5_3_msg;
  wire [7:0] weight_inter_5_4_msg;
  wire [7:0] weight_inter_5_5_msg;
  wire [7:0] weight_inter_5_6_msg;
  wire [7:0] weight_inter_5_7_msg;
  wire [7:0] weight_inter_6_0_msg;
  wire [7:0] weight_inter_6_1_msg;
  wire [7:0] weight_inter_6_2_msg;
  wire [7:0] weight_inter_6_3_msg;
  wire [7:0] weight_inter_6_4_msg;
  wire [7:0] weight_inter_6_5_msg;
  wire [7:0] weight_inter_6_6_msg;
  wire [7:0] weight_inter_6_7_msg;
  wire [7:0] weight_inter_7_0_msg;
  wire [7:0] weight_inter_7_1_msg;
  wire [7:0] weight_inter_7_2_msg;
  wire [7:0] weight_inter_7_3_msg;
  wire [7:0] weight_inter_7_4_msg;
  wire [7:0] weight_inter_7_5_msg;
  wire [7:0] weight_inter_7_6_msg;
  wire [7:0] weight_inter_7_7_msg;
  wire act_inter_0_0_val;
  wire act_inter_0_1_val;
  wire act_inter_0_2_val;
  wire act_inter_0_3_val;
  wire act_inter_0_4_val;
  wire act_inter_0_5_val;
  wire act_inter_0_6_val;
  wire act_inter_0_7_val;
  wire act_inter_1_0_val;
  wire act_inter_1_1_val;
  wire act_inter_1_2_val;
  wire act_inter_1_3_val;
  wire act_inter_1_4_val;
  wire act_inter_1_5_val;
  wire act_inter_1_6_val;
  wire act_inter_1_7_val;
  wire act_inter_2_0_val;
  wire act_inter_2_1_val;
  wire act_inter_2_2_val;
  wire act_inter_2_3_val;
  wire act_inter_2_4_val;
  wire act_inter_2_5_val;
  wire act_inter_2_6_val;
  wire act_inter_2_7_val;
  wire act_inter_3_0_val;
  wire act_inter_3_1_val;
  wire act_inter_3_2_val;
  wire act_inter_3_3_val;
  wire act_inter_3_4_val;
  wire act_inter_3_5_val;
  wire act_inter_3_6_val;
  wire act_inter_3_7_val;
  wire act_inter_4_0_val;
  wire act_inter_4_1_val;
  wire act_inter_4_2_val;
  wire act_inter_4_3_val;
  wire act_inter_4_4_val;
  wire act_inter_4_5_val;
  wire act_inter_4_6_val;
  wire act_inter_4_7_val;
  wire act_inter_5_0_val;
  wire act_inter_5_1_val;
  wire act_inter_5_2_val;
  wire act_inter_5_3_val;
  wire act_inter_5_4_val;
  wire act_inter_5_5_val;
  wire act_inter_5_6_val;
  wire act_inter_5_7_val;
  wire act_inter_6_0_val;
  wire act_inter_6_1_val;
  wire act_inter_6_2_val;
  wire act_inter_6_3_val;
  wire act_inter_6_4_val;
  wire act_inter_6_5_val;
  wire act_inter_6_6_val;
  wire act_inter_6_7_val;
  wire act_inter_7_0_val;
  wire act_inter_7_1_val;
  wire act_inter_7_2_val;
  wire act_inter_7_3_val;
  wire act_inter_7_4_val;
  wire act_inter_7_5_val;
  wire act_inter_7_6_val;
  wire act_inter_7_7_val;
  wire act_inter_0_0_rdy;
  wire act_inter_0_1_rdy;
  wire act_inter_0_2_rdy;
  wire act_inter_0_3_rdy;
  wire act_inter_0_4_rdy;
  wire act_inter_0_5_rdy;
  wire act_inter_0_6_rdy;
  wire act_inter_0_7_rdy;
  wire act_inter_1_0_rdy;
  wire act_inter_1_1_rdy;
  wire act_inter_1_2_rdy;
  wire act_inter_1_3_rdy;
  wire act_inter_1_4_rdy;
  wire act_inter_1_5_rdy;
  wire act_inter_1_6_rdy;
  wire act_inter_1_7_rdy;
  wire act_inter_2_0_rdy;
  wire act_inter_2_1_rdy;
  wire act_inter_2_2_rdy;
  wire act_inter_2_3_rdy;
  wire act_inter_2_4_rdy;
  wire act_inter_2_5_rdy;
  wire act_inter_2_6_rdy;
  wire act_inter_2_7_rdy;
  wire act_inter_3_0_rdy;
  wire act_inter_3_1_rdy;
  wire act_inter_3_2_rdy;
  wire act_inter_3_3_rdy;
  wire act_inter_3_4_rdy;
  wire act_inter_3_5_rdy;
  wire act_inter_3_6_rdy;
  wire act_inter_3_7_rdy;
  wire act_inter_4_0_rdy;
  wire act_inter_4_1_rdy;
  wire act_inter_4_2_rdy;
  wire act_inter_4_3_rdy;
  wire act_inter_4_4_rdy;
  wire act_inter_4_5_rdy;
  wire act_inter_4_6_rdy;
  wire act_inter_4_7_rdy;
  wire act_inter_5_0_rdy;
  wire act_inter_5_1_rdy;
  wire act_inter_5_2_rdy;
  wire act_inter_5_3_rdy;
  wire act_inter_5_4_rdy;
  wire act_inter_5_5_rdy;
  wire act_inter_5_6_rdy;
  wire act_inter_5_7_rdy;
  wire act_inter_6_0_rdy;
  wire act_inter_6_1_rdy;
  wire act_inter_6_2_rdy;
  wire act_inter_6_3_rdy;
  wire act_inter_6_4_rdy;
  wire act_inter_6_5_rdy;
  wire act_inter_6_6_rdy;
  wire act_inter_6_7_rdy;
  wire act_inter_7_0_rdy;
  wire act_inter_7_1_rdy;
  wire act_inter_7_2_rdy;
  wire act_inter_7_3_rdy;
  wire act_inter_7_4_rdy;
  wire act_inter_7_5_rdy;
  wire act_inter_7_6_rdy;
  wire act_inter_7_7_rdy;
  wire [7:0] act_inter_0_0_msg;
  wire [7:0] act_inter_0_1_msg;
  wire [7:0] act_inter_0_2_msg;
  wire [7:0] act_inter_0_3_msg;
  wire [7:0] act_inter_0_4_msg;
  wire [7:0] act_inter_0_5_msg;
  wire [7:0] act_inter_0_6_msg;
  wire [7:0] act_inter_0_7_msg;
  wire [7:0] act_inter_1_0_msg;
  wire [7:0] act_inter_1_1_msg;
  wire [7:0] act_inter_1_2_msg;
  wire [7:0] act_inter_1_3_msg;
  wire [7:0] act_inter_1_4_msg;
  wire [7:0] act_inter_1_5_msg;
  wire [7:0] act_inter_1_6_msg;
  wire [7:0] act_inter_1_7_msg;
  wire [7:0] act_inter_2_0_msg;
  wire [7:0] act_inter_2_1_msg;
  wire [7:0] act_inter_2_2_msg;
  wire [7:0] act_inter_2_3_msg;
  wire [7:0] act_inter_2_4_msg;
  wire [7:0] act_inter_2_5_msg;
  wire [7:0] act_inter_2_6_msg;
  wire [7:0] act_inter_2_7_msg;
  wire [7:0] act_inter_3_0_msg;
  wire [7:0] act_inter_3_1_msg;
  wire [7:0] act_inter_3_2_msg;
  wire [7:0] act_inter_3_3_msg;
  wire [7:0] act_inter_3_4_msg;
  wire [7:0] act_inter_3_5_msg;
  wire [7:0] act_inter_3_6_msg;
  wire [7:0] act_inter_3_7_msg;
  wire [7:0] act_inter_4_0_msg;
  wire [7:0] act_inter_4_1_msg;
  wire [7:0] act_inter_4_2_msg;
  wire [7:0] act_inter_4_3_msg;
  wire [7:0] act_inter_4_4_msg;
  wire [7:0] act_inter_4_5_msg;
  wire [7:0] act_inter_4_6_msg;
  wire [7:0] act_inter_4_7_msg;
  wire [7:0] act_inter_5_0_msg;
  wire [7:0] act_inter_5_1_msg;
  wire [7:0] act_inter_5_2_msg;
  wire [7:0] act_inter_5_3_msg;
  wire [7:0] act_inter_5_4_msg;
  wire [7:0] act_inter_5_5_msg;
  wire [7:0] act_inter_5_6_msg;
  wire [7:0] act_inter_5_7_msg;
  wire [7:0] act_inter_6_0_msg;
  wire [7:0] act_inter_6_1_msg;
  wire [7:0] act_inter_6_2_msg;
  wire [7:0] act_inter_6_3_msg;
  wire [7:0] act_inter_6_4_msg;
  wire [7:0] act_inter_6_5_msg;
  wire [7:0] act_inter_6_6_msg;
  wire [7:0] act_inter_6_7_msg;
  wire [7:0] act_inter_7_0_msg;
  wire [7:0] act_inter_7_1_msg;
  wire [7:0] act_inter_7_2_msg;
  wire [7:0] act_inter_7_3_msg;
  wire [7:0] act_inter_7_4_msg;
  wire [7:0] act_inter_7_5_msg;
  wire [7:0] act_inter_7_6_msg;
  wire [7:0] act_inter_7_7_msg;
  wire accum_inter_0_0_val;
  wire accum_inter_0_1_val;
  wire accum_inter_0_2_val;
  wire accum_inter_0_3_val;
  wire accum_inter_0_4_val;
  wire accum_inter_0_5_val;
  wire accum_inter_0_6_val;
  wire accum_inter_0_7_val;
  wire accum_inter_1_0_val;
  wire accum_inter_1_1_val;
  wire accum_inter_1_2_val;
  wire accum_inter_1_3_val;
  wire accum_inter_1_4_val;
  wire accum_inter_1_5_val;
  wire accum_inter_1_6_val;
  wire accum_inter_1_7_val;
  wire accum_inter_2_0_val;
  wire accum_inter_2_1_val;
  wire accum_inter_2_2_val;
  wire accum_inter_2_3_val;
  wire accum_inter_2_4_val;
  wire accum_inter_2_5_val;
  wire accum_inter_2_6_val;
  wire accum_inter_2_7_val;
  wire accum_inter_3_0_val;
  wire accum_inter_3_1_val;
  wire accum_inter_3_2_val;
  wire accum_inter_3_3_val;
  wire accum_inter_3_4_val;
  wire accum_inter_3_5_val;
  wire accum_inter_3_6_val;
  wire accum_inter_3_7_val;
  wire accum_inter_4_0_val;
  wire accum_inter_4_1_val;
  wire accum_inter_4_2_val;
  wire accum_inter_4_3_val;
  wire accum_inter_4_4_val;
  wire accum_inter_4_5_val;
  wire accum_inter_4_6_val;
  wire accum_inter_4_7_val;
  wire accum_inter_5_0_val;
  wire accum_inter_5_1_val;
  wire accum_inter_5_2_val;
  wire accum_inter_5_3_val;
  wire accum_inter_5_4_val;
  wire accum_inter_5_5_val;
  wire accum_inter_5_6_val;
  wire accum_inter_5_7_val;
  wire accum_inter_6_0_val;
  wire accum_inter_6_1_val;
  wire accum_inter_6_2_val;
  wire accum_inter_6_3_val;
  wire accum_inter_6_4_val;
  wire accum_inter_6_5_val;
  wire accum_inter_6_6_val;
  wire accum_inter_6_7_val;
  wire accum_inter_7_0_val;
  wire accum_inter_7_1_val;
  wire accum_inter_7_2_val;
  wire accum_inter_7_3_val;
  wire accum_inter_7_4_val;
  wire accum_inter_7_5_val;
  wire accum_inter_7_6_val;
  wire accum_inter_7_7_val;
  wire accum_inter_0_0_rdy;
  wire accum_inter_0_1_rdy;
  wire accum_inter_0_2_rdy;
  wire accum_inter_0_3_rdy;
  wire accum_inter_0_4_rdy;
  wire accum_inter_0_5_rdy;
  wire accum_inter_0_6_rdy;
  wire accum_inter_0_7_rdy;
  wire accum_inter_1_0_rdy;
  wire accum_inter_1_1_rdy;
  wire accum_inter_1_2_rdy;
  wire accum_inter_1_3_rdy;
  wire accum_inter_1_4_rdy;
  wire accum_inter_1_5_rdy;
  wire accum_inter_1_6_rdy;
  wire accum_inter_1_7_rdy;
  wire accum_inter_2_0_rdy;
  wire accum_inter_2_1_rdy;
  wire accum_inter_2_2_rdy;
  wire accum_inter_2_3_rdy;
  wire accum_inter_2_4_rdy;
  wire accum_inter_2_5_rdy;
  wire accum_inter_2_6_rdy;
  wire accum_inter_2_7_rdy;
  wire accum_inter_3_0_rdy;
  wire accum_inter_3_1_rdy;
  wire accum_inter_3_2_rdy;
  wire accum_inter_3_3_rdy;
  wire accum_inter_3_4_rdy;
  wire accum_inter_3_5_rdy;
  wire accum_inter_3_6_rdy;
  wire accum_inter_3_7_rdy;
  wire accum_inter_4_0_rdy;
  wire accum_inter_4_1_rdy;
  wire accum_inter_4_2_rdy;
  wire accum_inter_4_3_rdy;
  wire accum_inter_4_4_rdy;
  wire accum_inter_4_5_rdy;
  wire accum_inter_4_6_rdy;
  wire accum_inter_4_7_rdy;
  wire accum_inter_5_0_rdy;
  wire accum_inter_5_1_rdy;
  wire accum_inter_5_2_rdy;
  wire accum_inter_5_3_rdy;
  wire accum_inter_5_4_rdy;
  wire accum_inter_5_5_rdy;
  wire accum_inter_5_6_rdy;
  wire accum_inter_5_7_rdy;
  wire accum_inter_6_0_rdy;
  wire accum_inter_6_1_rdy;
  wire accum_inter_6_2_rdy;
  wire accum_inter_6_3_rdy;
  wire accum_inter_6_4_rdy;
  wire accum_inter_6_5_rdy;
  wire accum_inter_6_6_rdy;
  wire accum_inter_6_7_rdy;
  wire accum_inter_7_0_rdy;
  wire accum_inter_7_1_rdy;
  wire accum_inter_7_2_rdy;
  wire accum_inter_7_3_rdy;
  wire accum_inter_7_4_rdy;
  wire accum_inter_7_5_rdy;
  wire accum_inter_7_6_rdy;
  wire accum_inter_7_7_rdy;
  wire [31:0] accum_inter_0_0_msg;
  wire [31:0] accum_inter_0_1_msg;
  wire [31:0] accum_inter_0_2_msg;
  wire [31:0] accum_inter_0_3_msg;
  wire [31:0] accum_inter_0_4_msg;
  wire [31:0] accum_inter_0_5_msg;
  wire [31:0] accum_inter_0_6_msg;
  wire [31:0] accum_inter_0_7_msg;
  wire [31:0] accum_inter_1_0_msg;
  wire [31:0] accum_inter_1_1_msg;
  wire [31:0] accum_inter_1_2_msg;
  wire [31:0] accum_inter_1_3_msg;
  wire [31:0] accum_inter_1_4_msg;
  wire [31:0] accum_inter_1_5_msg;
  wire [31:0] accum_inter_1_6_msg;
  wire [31:0] accum_inter_1_7_msg;
  wire [31:0] accum_inter_2_0_msg;
  wire [31:0] accum_inter_2_1_msg;
  wire [31:0] accum_inter_2_2_msg;
  wire [31:0] accum_inter_2_3_msg;
  wire [31:0] accum_inter_2_4_msg;
  wire [31:0] accum_inter_2_5_msg;
  wire [31:0] accum_inter_2_6_msg;
  wire [31:0] accum_inter_2_7_msg;
  wire [31:0] accum_inter_3_0_msg;
  wire [31:0] accum_inter_3_1_msg;
  wire [31:0] accum_inter_3_2_msg;
  wire [31:0] accum_inter_3_3_msg;
  wire [31:0] accum_inter_3_4_msg;
  wire [31:0] accum_inter_3_5_msg;
  wire [31:0] accum_inter_3_6_msg;
  wire [31:0] accum_inter_3_7_msg;
  wire [31:0] accum_inter_4_0_msg;
  wire [31:0] accum_inter_4_1_msg;
  wire [31:0] accum_inter_4_2_msg;
  wire [31:0] accum_inter_4_3_msg;
  wire [31:0] accum_inter_4_4_msg;
  wire [31:0] accum_inter_4_5_msg;
  wire [31:0] accum_inter_4_6_msg;
  wire [31:0] accum_inter_4_7_msg;
  wire [31:0] accum_inter_5_0_msg;
  wire [31:0] accum_inter_5_1_msg;
  wire [31:0] accum_inter_5_2_msg;
  wire [31:0] accum_inter_5_3_msg;
  wire [31:0] accum_inter_5_4_msg;
  wire [31:0] accum_inter_5_5_msg;
  wire [31:0] accum_inter_5_6_msg;
  wire [31:0] accum_inter_5_7_msg;
  wire [31:0] accum_inter_6_0_msg;
  wire [31:0] accum_inter_6_1_msg;
  wire [31:0] accum_inter_6_2_msg;
  wire [31:0] accum_inter_6_3_msg;
  wire [31:0] accum_inter_6_4_msg;
  wire [31:0] accum_inter_6_5_msg;
  wire [31:0] accum_inter_6_6_msg;
  wire [31:0] accum_inter_6_7_msg;
  wire [31:0] accum_inter_7_0_msg;
  wire [31:0] accum_inter_7_1_msg;
  wire [31:0] accum_inter_7_2_msg;
  wire [31:0] accum_inter_7_3_msg;
  wire [31:0] accum_inter_7_4_msg;
  wire [31:0] accum_inter_7_5_msg;
  wire [31:0] accum_inter_7_6_msg;
  wire [31:0] accum_inter_7_7_msg;
  wire [7:0] act_inter_PopNB_7_mioi_data_rsc_z;
  wire act_inter_PopNB_7_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_15_mioi_data_rsc_z;
  wire act_inter_PopNB_15_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_23_mioi_data_rsc_z;
  wire act_inter_PopNB_23_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_31_mioi_data_rsc_z;
  wire act_inter_PopNB_31_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_39_mioi_data_rsc_z;
  wire act_inter_PopNB_39_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_47_mioi_data_rsc_z;
  wire act_inter_PopNB_47_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_55_mioi_data_rsc_z;
  wire act_inter_PopNB_55_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_63_mioi_data_rsc_z;
  wire act_inter_PopNB_63_mioi_return_rsc_z;
  wire accum_inter_PushNB_mioi_return_rsc_z;
  wire accum_inter_PushNB_1_mioi_return_rsc_z;
  wire accum_inter_PushNB_2_mioi_return_rsc_z;
  wire accum_inter_PushNB_3_mioi_return_rsc_z;
  wire accum_inter_PushNB_4_mioi_return_rsc_z;
  wire accum_inter_PushNB_5_mioi_return_rsc_z;
  wire accum_inter_PushNB_6_mioi_return_rsc_z;
  wire accum_inter_PushNB_7_mioi_return_rsc_z;
  wire act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff;
  wire accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_7_mioi
      (
      .this_val(act_inter_0_7_val),
      .this_rdy(act_inter_0_7_rdy),
      .this_msg(act_inter_0_7_msg),
      .data_rsc_z(act_inter_PopNB_7_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_7_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_15_mioi
      (
      .this_val(act_inter_1_7_val),
      .this_rdy(act_inter_1_7_rdy),
      .this_msg(act_inter_1_7_msg),
      .data_rsc_z(act_inter_PopNB_15_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_15_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_23_mioi
      (
      .this_val(act_inter_2_7_val),
      .this_rdy(act_inter_2_7_rdy),
      .this_msg(act_inter_2_7_msg),
      .data_rsc_z(act_inter_PopNB_23_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_23_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_31_mioi
      (
      .this_val(act_inter_3_7_val),
      .this_rdy(act_inter_3_7_rdy),
      .this_msg(act_inter_3_7_msg),
      .data_rsc_z(act_inter_PopNB_31_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_31_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_39_mioi
      (
      .this_val(act_inter_4_7_val),
      .this_rdy(act_inter_4_7_rdy),
      .this_msg(act_inter_4_7_msg),
      .data_rsc_z(act_inter_PopNB_39_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_39_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_47_mioi
      (
      .this_val(act_inter_5_7_val),
      .this_rdy(act_inter_5_7_rdy),
      .this_msg(act_inter_5_7_msg),
      .data_rsc_z(act_inter_PopNB_47_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_47_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_55_mioi
      (
      .this_val(act_inter_6_7_val),
      .this_rdy(act_inter_6_7_rdy),
      .this_msg(act_inter_6_7_msg),
      .data_rsc_z(act_inter_PopNB_55_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_55_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_63_mioi
      (
      .this_val(act_inter_7_7_val),
      .this_rdy(act_inter_7_7_rdy),
      .this_msg(act_inter_7_7_msg),
      .data_rsc_z(act_inter_PopNB_63_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_63_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_mioi
      (
      .this_val(accum_inter_0_0_val),
      .this_rdy(accum_inter_0_0_rdy),
      .this_msg(accum_inter_0_0_msg),
      .return_rsc_z(accum_inter_PushNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_1_mioi
      (
      .this_val(accum_inter_0_1_val),
      .this_rdy(accum_inter_0_1_rdy),
      .this_msg(accum_inter_0_1_msg),
      .return_rsc_z(accum_inter_PushNB_1_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_2_mioi
      (
      .this_val(accum_inter_0_2_val),
      .this_rdy(accum_inter_0_2_rdy),
      .this_msg(accum_inter_0_2_msg),
      .return_rsc_z(accum_inter_PushNB_2_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_3_mioi
      (
      .this_val(accum_inter_0_3_val),
      .this_rdy(accum_inter_0_3_rdy),
      .this_msg(accum_inter_0_3_msg),
      .return_rsc_z(accum_inter_PushNB_3_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_4_mioi
      (
      .this_val(accum_inter_0_4_val),
      .this_rdy(accum_inter_0_4_rdy),
      .this_msg(accum_inter_0_4_msg),
      .return_rsc_z(accum_inter_PushNB_4_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_5_mioi
      (
      .this_val(accum_inter_0_5_val),
      .this_rdy(accum_inter_0_5_rdy),
      .this_msg(accum_inter_0_5_msg),
      .return_rsc_z(accum_inter_PushNB_5_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_6_mioi
      (
      .this_val(accum_inter_0_6_val),
      .this_rdy(accum_inter_0_6_rdy),
      .this_msg(accum_inter_0_6_msg),
      .return_rsc_z(accum_inter_PushNB_6_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_7_mioi
      (
      .this_val(accum_inter_0_7_val),
      .this_rdy(accum_inter_0_7_rdy),
      .this_msg(accum_inter_0_7_msg),
      .return_rsc_z(accum_inter_PushNB_7_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  SysPE SysPE_1 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_0_val),
      .weight_in_rdy(weight_in_vec_0_rdy),
      .weight_in_msg(weight_in_vec_0_msg),
      .act_in_val(act_in_vec_0_val),
      .act_in_rdy(act_in_vec_0_rdy),
      .act_in_msg(act_in_vec_0_msg),
      .accum_in_val(accum_inter_0_0_val),
      .accum_in_rdy(accum_inter_0_0_rdy),
      .accum_in_msg(accum_inter_0_0_msg),
      .weight_out_val(weight_inter_0_0_val),
      .weight_out_rdy(weight_inter_0_0_rdy),
      .weight_out_msg(weight_inter_0_0_msg),
      .act_out_val(act_inter_0_0_val),
      .act_out_rdy(act_inter_0_0_rdy),
      .act_out_msg(act_inter_0_0_msg),
      .accum_out_val(accum_inter_1_0_val),
      .accum_out_rdy(accum_inter_1_0_rdy),
      .accum_out_msg(accum_inter_1_0_msg)
    );
  SysPE SysPE_2 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_1_val),
      .weight_in_rdy(weight_in_vec_1_rdy),
      .weight_in_msg(weight_in_vec_1_msg),
      .act_in_val(act_inter_0_0_val),
      .act_in_rdy(act_inter_0_0_rdy),
      .act_in_msg(act_inter_0_0_msg),
      .accum_in_val(accum_inter_0_1_val),
      .accum_in_rdy(accum_inter_0_1_rdy),
      .accum_in_msg(accum_inter_0_1_msg),
      .weight_out_val(weight_inter_0_1_val),
      .weight_out_rdy(weight_inter_0_1_rdy),
      .weight_out_msg(weight_inter_0_1_msg),
      .act_out_val(act_inter_0_1_val),
      .act_out_rdy(act_inter_0_1_rdy),
      .act_out_msg(act_inter_0_1_msg),
      .accum_out_val(accum_inter_1_1_val),
      .accum_out_rdy(accum_inter_1_1_rdy),
      .accum_out_msg(accum_inter_1_1_msg)
    );
  SysPE SysPE_3 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_2_val),
      .weight_in_rdy(weight_in_vec_2_rdy),
      .weight_in_msg(weight_in_vec_2_msg),
      .act_in_val(act_inter_0_1_val),
      .act_in_rdy(act_inter_0_1_rdy),
      .act_in_msg(act_inter_0_1_msg),
      .accum_in_val(accum_inter_0_2_val),
      .accum_in_rdy(accum_inter_0_2_rdy),
      .accum_in_msg(accum_inter_0_2_msg),
      .weight_out_val(weight_inter_0_2_val),
      .weight_out_rdy(weight_inter_0_2_rdy),
      .weight_out_msg(weight_inter_0_2_msg),
      .act_out_val(act_inter_0_2_val),
      .act_out_rdy(act_inter_0_2_rdy),
      .act_out_msg(act_inter_0_2_msg),
      .accum_out_val(accum_inter_1_2_val),
      .accum_out_rdy(accum_inter_1_2_rdy),
      .accum_out_msg(accum_inter_1_2_msg)
    );
  SysPE SysPE_4 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_3_val),
      .weight_in_rdy(weight_in_vec_3_rdy),
      .weight_in_msg(weight_in_vec_3_msg),
      .act_in_val(act_inter_0_2_val),
      .act_in_rdy(act_inter_0_2_rdy),
      .act_in_msg(act_inter_0_2_msg),
      .accum_in_val(accum_inter_0_3_val),
      .accum_in_rdy(accum_inter_0_3_rdy),
      .accum_in_msg(accum_inter_0_3_msg),
      .weight_out_val(weight_inter_0_3_val),
      .weight_out_rdy(weight_inter_0_3_rdy),
      .weight_out_msg(weight_inter_0_3_msg),
      .act_out_val(act_inter_0_3_val),
      .act_out_rdy(act_inter_0_3_rdy),
      .act_out_msg(act_inter_0_3_msg),
      .accum_out_val(accum_inter_1_3_val),
      .accum_out_rdy(accum_inter_1_3_rdy),
      .accum_out_msg(accum_inter_1_3_msg)
    );
  SysPE SysPE_5 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_4_val),
      .weight_in_rdy(weight_in_vec_4_rdy),
      .weight_in_msg(weight_in_vec_4_msg),
      .act_in_val(act_inter_0_3_val),
      .act_in_rdy(act_inter_0_3_rdy),
      .act_in_msg(act_inter_0_3_msg),
      .accum_in_val(accum_inter_0_4_val),
      .accum_in_rdy(accum_inter_0_4_rdy),
      .accum_in_msg(accum_inter_0_4_msg),
      .weight_out_val(weight_inter_0_4_val),
      .weight_out_rdy(weight_inter_0_4_rdy),
      .weight_out_msg(weight_inter_0_4_msg),
      .act_out_val(act_inter_0_4_val),
      .act_out_rdy(act_inter_0_4_rdy),
      .act_out_msg(act_inter_0_4_msg),
      .accum_out_val(accum_inter_1_4_val),
      .accum_out_rdy(accum_inter_1_4_rdy),
      .accum_out_msg(accum_inter_1_4_msg)
    );
  SysPE SysPE_6 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_5_val),
      .weight_in_rdy(weight_in_vec_5_rdy),
      .weight_in_msg(weight_in_vec_5_msg),
      .act_in_val(act_inter_0_4_val),
      .act_in_rdy(act_inter_0_4_rdy),
      .act_in_msg(act_inter_0_4_msg),
      .accum_in_val(accum_inter_0_5_val),
      .accum_in_rdy(accum_inter_0_5_rdy),
      .accum_in_msg(accum_inter_0_5_msg),
      .weight_out_val(weight_inter_0_5_val),
      .weight_out_rdy(weight_inter_0_5_rdy),
      .weight_out_msg(weight_inter_0_5_msg),
      .act_out_val(act_inter_0_5_val),
      .act_out_rdy(act_inter_0_5_rdy),
      .act_out_msg(act_inter_0_5_msg),
      .accum_out_val(accum_inter_1_5_val),
      .accum_out_rdy(accum_inter_1_5_rdy),
      .accum_out_msg(accum_inter_1_5_msg)
    );
  SysPE SysPE_7 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_6_val),
      .weight_in_rdy(weight_in_vec_6_rdy),
      .weight_in_msg(weight_in_vec_6_msg),
      .act_in_val(act_inter_0_5_val),
      .act_in_rdy(act_inter_0_5_rdy),
      .act_in_msg(act_inter_0_5_msg),
      .accum_in_val(accum_inter_0_6_val),
      .accum_in_rdy(accum_inter_0_6_rdy),
      .accum_in_msg(accum_inter_0_6_msg),
      .weight_out_val(weight_inter_0_6_val),
      .weight_out_rdy(weight_inter_0_6_rdy),
      .weight_out_msg(weight_inter_0_6_msg),
      .act_out_val(act_inter_0_6_val),
      .act_out_rdy(act_inter_0_6_rdy),
      .act_out_msg(act_inter_0_6_msg),
      .accum_out_val(accum_inter_1_6_val),
      .accum_out_rdy(accum_inter_1_6_rdy),
      .accum_out_msg(accum_inter_1_6_msg)
    );
  SysPE SysPE_8 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_7_val),
      .weight_in_rdy(weight_in_vec_7_rdy),
      .weight_in_msg(weight_in_vec_7_msg),
      .act_in_val(act_inter_0_6_val),
      .act_in_rdy(act_inter_0_6_rdy),
      .act_in_msg(act_inter_0_6_msg),
      .accum_in_val(accum_inter_0_7_val),
      .accum_in_rdy(accum_inter_0_7_rdy),
      .accum_in_msg(accum_inter_0_7_msg),
      .weight_out_val(weight_inter_0_7_val),
      .weight_out_rdy(weight_inter_0_7_rdy),
      .weight_out_msg(weight_inter_0_7_msg),
      .act_out_val(act_inter_0_7_val),
      .act_out_rdy(act_inter_0_7_rdy),
      .act_out_msg(act_inter_0_7_msg),
      .accum_out_val(accum_inter_1_7_val),
      .accum_out_rdy(accum_inter_1_7_rdy),
      .accum_out_msg(accum_inter_1_7_msg)
    );
  SysPE SysPE_9 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_0_val),
      .weight_in_rdy(weight_inter_0_0_rdy),
      .weight_in_msg(weight_inter_0_0_msg),
      .act_in_val(act_in_vec_1_val),
      .act_in_rdy(act_in_vec_1_rdy),
      .act_in_msg(act_in_vec_1_msg),
      .accum_in_val(accum_inter_1_0_val),
      .accum_in_rdy(accum_inter_1_0_rdy),
      .accum_in_msg(accum_inter_1_0_msg),
      .weight_out_val(weight_inter_1_0_val),
      .weight_out_rdy(weight_inter_1_0_rdy),
      .weight_out_msg(weight_inter_1_0_msg),
      .act_out_val(act_inter_1_0_val),
      .act_out_rdy(act_inter_1_0_rdy),
      .act_out_msg(act_inter_1_0_msg),
      .accum_out_val(accum_inter_2_0_val),
      .accum_out_rdy(accum_inter_2_0_rdy),
      .accum_out_msg(accum_inter_2_0_msg)
    );
  SysPE SysPE_10 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_1_val),
      .weight_in_rdy(weight_inter_0_1_rdy),
      .weight_in_msg(weight_inter_0_1_msg),
      .act_in_val(act_inter_1_0_val),
      .act_in_rdy(act_inter_1_0_rdy),
      .act_in_msg(act_inter_1_0_msg),
      .accum_in_val(accum_inter_1_1_val),
      .accum_in_rdy(accum_inter_1_1_rdy),
      .accum_in_msg(accum_inter_1_1_msg),
      .weight_out_val(weight_inter_1_1_val),
      .weight_out_rdy(weight_inter_1_1_rdy),
      .weight_out_msg(weight_inter_1_1_msg),
      .act_out_val(act_inter_1_1_val),
      .act_out_rdy(act_inter_1_1_rdy),
      .act_out_msg(act_inter_1_1_msg),
      .accum_out_val(accum_inter_2_1_val),
      .accum_out_rdy(accum_inter_2_1_rdy),
      .accum_out_msg(accum_inter_2_1_msg)
    );
  SysPE SysPE_11 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_2_val),
      .weight_in_rdy(weight_inter_0_2_rdy),
      .weight_in_msg(weight_inter_0_2_msg),
      .act_in_val(act_inter_1_1_val),
      .act_in_rdy(act_inter_1_1_rdy),
      .act_in_msg(act_inter_1_1_msg),
      .accum_in_val(accum_inter_1_2_val),
      .accum_in_rdy(accum_inter_1_2_rdy),
      .accum_in_msg(accum_inter_1_2_msg),
      .weight_out_val(weight_inter_1_2_val),
      .weight_out_rdy(weight_inter_1_2_rdy),
      .weight_out_msg(weight_inter_1_2_msg),
      .act_out_val(act_inter_1_2_val),
      .act_out_rdy(act_inter_1_2_rdy),
      .act_out_msg(act_inter_1_2_msg),
      .accum_out_val(accum_inter_2_2_val),
      .accum_out_rdy(accum_inter_2_2_rdy),
      .accum_out_msg(accum_inter_2_2_msg)
    );
  SysPE SysPE_12 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_3_val),
      .weight_in_rdy(weight_inter_0_3_rdy),
      .weight_in_msg(weight_inter_0_3_msg),
      .act_in_val(act_inter_1_2_val),
      .act_in_rdy(act_inter_1_2_rdy),
      .act_in_msg(act_inter_1_2_msg),
      .accum_in_val(accum_inter_1_3_val),
      .accum_in_rdy(accum_inter_1_3_rdy),
      .accum_in_msg(accum_inter_1_3_msg),
      .weight_out_val(weight_inter_1_3_val),
      .weight_out_rdy(weight_inter_1_3_rdy),
      .weight_out_msg(weight_inter_1_3_msg),
      .act_out_val(act_inter_1_3_val),
      .act_out_rdy(act_inter_1_3_rdy),
      .act_out_msg(act_inter_1_3_msg),
      .accum_out_val(accum_inter_2_3_val),
      .accum_out_rdy(accum_inter_2_3_rdy),
      .accum_out_msg(accum_inter_2_3_msg)
    );
  SysPE SysPE_13 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_4_val),
      .weight_in_rdy(weight_inter_0_4_rdy),
      .weight_in_msg(weight_inter_0_4_msg),
      .act_in_val(act_inter_1_3_val),
      .act_in_rdy(act_inter_1_3_rdy),
      .act_in_msg(act_inter_1_3_msg),
      .accum_in_val(accum_inter_1_4_val),
      .accum_in_rdy(accum_inter_1_4_rdy),
      .accum_in_msg(accum_inter_1_4_msg),
      .weight_out_val(weight_inter_1_4_val),
      .weight_out_rdy(weight_inter_1_4_rdy),
      .weight_out_msg(weight_inter_1_4_msg),
      .act_out_val(act_inter_1_4_val),
      .act_out_rdy(act_inter_1_4_rdy),
      .act_out_msg(act_inter_1_4_msg),
      .accum_out_val(accum_inter_2_4_val),
      .accum_out_rdy(accum_inter_2_4_rdy),
      .accum_out_msg(accum_inter_2_4_msg)
    );
  SysPE SysPE_14 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_5_val),
      .weight_in_rdy(weight_inter_0_5_rdy),
      .weight_in_msg(weight_inter_0_5_msg),
      .act_in_val(act_inter_1_4_val),
      .act_in_rdy(act_inter_1_4_rdy),
      .act_in_msg(act_inter_1_4_msg),
      .accum_in_val(accum_inter_1_5_val),
      .accum_in_rdy(accum_inter_1_5_rdy),
      .accum_in_msg(accum_inter_1_5_msg),
      .weight_out_val(weight_inter_1_5_val),
      .weight_out_rdy(weight_inter_1_5_rdy),
      .weight_out_msg(weight_inter_1_5_msg),
      .act_out_val(act_inter_1_5_val),
      .act_out_rdy(act_inter_1_5_rdy),
      .act_out_msg(act_inter_1_5_msg),
      .accum_out_val(accum_inter_2_5_val),
      .accum_out_rdy(accum_inter_2_5_rdy),
      .accum_out_msg(accum_inter_2_5_msg)
    );
  SysPE SysPE_15 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_6_val),
      .weight_in_rdy(weight_inter_0_6_rdy),
      .weight_in_msg(weight_inter_0_6_msg),
      .act_in_val(act_inter_1_5_val),
      .act_in_rdy(act_inter_1_5_rdy),
      .act_in_msg(act_inter_1_5_msg),
      .accum_in_val(accum_inter_1_6_val),
      .accum_in_rdy(accum_inter_1_6_rdy),
      .accum_in_msg(accum_inter_1_6_msg),
      .weight_out_val(weight_inter_1_6_val),
      .weight_out_rdy(weight_inter_1_6_rdy),
      .weight_out_msg(weight_inter_1_6_msg),
      .act_out_val(act_inter_1_6_val),
      .act_out_rdy(act_inter_1_6_rdy),
      .act_out_msg(act_inter_1_6_msg),
      .accum_out_val(accum_inter_2_6_val),
      .accum_out_rdy(accum_inter_2_6_rdy),
      .accum_out_msg(accum_inter_2_6_msg)
    );
  SysPE SysPE_16 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_7_val),
      .weight_in_rdy(weight_inter_0_7_rdy),
      .weight_in_msg(weight_inter_0_7_msg),
      .act_in_val(act_inter_1_6_val),
      .act_in_rdy(act_inter_1_6_rdy),
      .act_in_msg(act_inter_1_6_msg),
      .accum_in_val(accum_inter_1_7_val),
      .accum_in_rdy(accum_inter_1_7_rdy),
      .accum_in_msg(accum_inter_1_7_msg),
      .weight_out_val(weight_inter_1_7_val),
      .weight_out_rdy(weight_inter_1_7_rdy),
      .weight_out_msg(weight_inter_1_7_msg),
      .act_out_val(act_inter_1_7_val),
      .act_out_rdy(act_inter_1_7_rdy),
      .act_out_msg(act_inter_1_7_msg),
      .accum_out_val(accum_inter_2_7_val),
      .accum_out_rdy(accum_inter_2_7_rdy),
      .accum_out_msg(accum_inter_2_7_msg)
    );
  SysPE SysPE_17 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_0_val),
      .weight_in_rdy(weight_inter_1_0_rdy),
      .weight_in_msg(weight_inter_1_0_msg),
      .act_in_val(act_in_vec_2_val),
      .act_in_rdy(act_in_vec_2_rdy),
      .act_in_msg(act_in_vec_2_msg),
      .accum_in_val(accum_inter_2_0_val),
      .accum_in_rdy(accum_inter_2_0_rdy),
      .accum_in_msg(accum_inter_2_0_msg),
      .weight_out_val(weight_inter_2_0_val),
      .weight_out_rdy(weight_inter_2_0_rdy),
      .weight_out_msg(weight_inter_2_0_msg),
      .act_out_val(act_inter_2_0_val),
      .act_out_rdy(act_inter_2_0_rdy),
      .act_out_msg(act_inter_2_0_msg),
      .accum_out_val(accum_inter_3_0_val),
      .accum_out_rdy(accum_inter_3_0_rdy),
      .accum_out_msg(accum_inter_3_0_msg)
    );
  SysPE SysPE_18 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_1_val),
      .weight_in_rdy(weight_inter_1_1_rdy),
      .weight_in_msg(weight_inter_1_1_msg),
      .act_in_val(act_inter_2_0_val),
      .act_in_rdy(act_inter_2_0_rdy),
      .act_in_msg(act_inter_2_0_msg),
      .accum_in_val(accum_inter_2_1_val),
      .accum_in_rdy(accum_inter_2_1_rdy),
      .accum_in_msg(accum_inter_2_1_msg),
      .weight_out_val(weight_inter_2_1_val),
      .weight_out_rdy(weight_inter_2_1_rdy),
      .weight_out_msg(weight_inter_2_1_msg),
      .act_out_val(act_inter_2_1_val),
      .act_out_rdy(act_inter_2_1_rdy),
      .act_out_msg(act_inter_2_1_msg),
      .accum_out_val(accum_inter_3_1_val),
      .accum_out_rdy(accum_inter_3_1_rdy),
      .accum_out_msg(accum_inter_3_1_msg)
    );
  SysPE SysPE_19 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_2_val),
      .weight_in_rdy(weight_inter_1_2_rdy),
      .weight_in_msg(weight_inter_1_2_msg),
      .act_in_val(act_inter_2_1_val),
      .act_in_rdy(act_inter_2_1_rdy),
      .act_in_msg(act_inter_2_1_msg),
      .accum_in_val(accum_inter_2_2_val),
      .accum_in_rdy(accum_inter_2_2_rdy),
      .accum_in_msg(accum_inter_2_2_msg),
      .weight_out_val(weight_inter_2_2_val),
      .weight_out_rdy(weight_inter_2_2_rdy),
      .weight_out_msg(weight_inter_2_2_msg),
      .act_out_val(act_inter_2_2_val),
      .act_out_rdy(act_inter_2_2_rdy),
      .act_out_msg(act_inter_2_2_msg),
      .accum_out_val(accum_inter_3_2_val),
      .accum_out_rdy(accum_inter_3_2_rdy),
      .accum_out_msg(accum_inter_3_2_msg)
    );
  SysPE SysPE_20 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_3_val),
      .weight_in_rdy(weight_inter_1_3_rdy),
      .weight_in_msg(weight_inter_1_3_msg),
      .act_in_val(act_inter_2_2_val),
      .act_in_rdy(act_inter_2_2_rdy),
      .act_in_msg(act_inter_2_2_msg),
      .accum_in_val(accum_inter_2_3_val),
      .accum_in_rdy(accum_inter_2_3_rdy),
      .accum_in_msg(accum_inter_2_3_msg),
      .weight_out_val(weight_inter_2_3_val),
      .weight_out_rdy(weight_inter_2_3_rdy),
      .weight_out_msg(weight_inter_2_3_msg),
      .act_out_val(act_inter_2_3_val),
      .act_out_rdy(act_inter_2_3_rdy),
      .act_out_msg(act_inter_2_3_msg),
      .accum_out_val(accum_inter_3_3_val),
      .accum_out_rdy(accum_inter_3_3_rdy),
      .accum_out_msg(accum_inter_3_3_msg)
    );
  SysPE SysPE_21 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_4_val),
      .weight_in_rdy(weight_inter_1_4_rdy),
      .weight_in_msg(weight_inter_1_4_msg),
      .act_in_val(act_inter_2_3_val),
      .act_in_rdy(act_inter_2_3_rdy),
      .act_in_msg(act_inter_2_3_msg),
      .accum_in_val(accum_inter_2_4_val),
      .accum_in_rdy(accum_inter_2_4_rdy),
      .accum_in_msg(accum_inter_2_4_msg),
      .weight_out_val(weight_inter_2_4_val),
      .weight_out_rdy(weight_inter_2_4_rdy),
      .weight_out_msg(weight_inter_2_4_msg),
      .act_out_val(act_inter_2_4_val),
      .act_out_rdy(act_inter_2_4_rdy),
      .act_out_msg(act_inter_2_4_msg),
      .accum_out_val(accum_inter_3_4_val),
      .accum_out_rdy(accum_inter_3_4_rdy),
      .accum_out_msg(accum_inter_3_4_msg)
    );
  SysPE SysPE_22 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_5_val),
      .weight_in_rdy(weight_inter_1_5_rdy),
      .weight_in_msg(weight_inter_1_5_msg),
      .act_in_val(act_inter_2_4_val),
      .act_in_rdy(act_inter_2_4_rdy),
      .act_in_msg(act_inter_2_4_msg),
      .accum_in_val(accum_inter_2_5_val),
      .accum_in_rdy(accum_inter_2_5_rdy),
      .accum_in_msg(accum_inter_2_5_msg),
      .weight_out_val(weight_inter_2_5_val),
      .weight_out_rdy(weight_inter_2_5_rdy),
      .weight_out_msg(weight_inter_2_5_msg),
      .act_out_val(act_inter_2_5_val),
      .act_out_rdy(act_inter_2_5_rdy),
      .act_out_msg(act_inter_2_5_msg),
      .accum_out_val(accum_inter_3_5_val),
      .accum_out_rdy(accum_inter_3_5_rdy),
      .accum_out_msg(accum_inter_3_5_msg)
    );
  SysPE SysPE_23 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_6_val),
      .weight_in_rdy(weight_inter_1_6_rdy),
      .weight_in_msg(weight_inter_1_6_msg),
      .act_in_val(act_inter_2_5_val),
      .act_in_rdy(act_inter_2_5_rdy),
      .act_in_msg(act_inter_2_5_msg),
      .accum_in_val(accum_inter_2_6_val),
      .accum_in_rdy(accum_inter_2_6_rdy),
      .accum_in_msg(accum_inter_2_6_msg),
      .weight_out_val(weight_inter_2_6_val),
      .weight_out_rdy(weight_inter_2_6_rdy),
      .weight_out_msg(weight_inter_2_6_msg),
      .act_out_val(act_inter_2_6_val),
      .act_out_rdy(act_inter_2_6_rdy),
      .act_out_msg(act_inter_2_6_msg),
      .accum_out_val(accum_inter_3_6_val),
      .accum_out_rdy(accum_inter_3_6_rdy),
      .accum_out_msg(accum_inter_3_6_msg)
    );
  SysPE SysPE_24 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_7_val),
      .weight_in_rdy(weight_inter_1_7_rdy),
      .weight_in_msg(weight_inter_1_7_msg),
      .act_in_val(act_inter_2_6_val),
      .act_in_rdy(act_inter_2_6_rdy),
      .act_in_msg(act_inter_2_6_msg),
      .accum_in_val(accum_inter_2_7_val),
      .accum_in_rdy(accum_inter_2_7_rdy),
      .accum_in_msg(accum_inter_2_7_msg),
      .weight_out_val(weight_inter_2_7_val),
      .weight_out_rdy(weight_inter_2_7_rdy),
      .weight_out_msg(weight_inter_2_7_msg),
      .act_out_val(act_inter_2_7_val),
      .act_out_rdy(act_inter_2_7_rdy),
      .act_out_msg(act_inter_2_7_msg),
      .accum_out_val(accum_inter_3_7_val),
      .accum_out_rdy(accum_inter_3_7_rdy),
      .accum_out_msg(accum_inter_3_7_msg)
    );
  SysPE SysPE_25 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_0_val),
      .weight_in_rdy(weight_inter_2_0_rdy),
      .weight_in_msg(weight_inter_2_0_msg),
      .act_in_val(act_in_vec_3_val),
      .act_in_rdy(act_in_vec_3_rdy),
      .act_in_msg(act_in_vec_3_msg),
      .accum_in_val(accum_inter_3_0_val),
      .accum_in_rdy(accum_inter_3_0_rdy),
      .accum_in_msg(accum_inter_3_0_msg),
      .weight_out_val(weight_inter_3_0_val),
      .weight_out_rdy(weight_inter_3_0_rdy),
      .weight_out_msg(weight_inter_3_0_msg),
      .act_out_val(act_inter_3_0_val),
      .act_out_rdy(act_inter_3_0_rdy),
      .act_out_msg(act_inter_3_0_msg),
      .accum_out_val(accum_inter_4_0_val),
      .accum_out_rdy(accum_inter_4_0_rdy),
      .accum_out_msg(accum_inter_4_0_msg)
    );
  SysPE SysPE_26 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_1_val),
      .weight_in_rdy(weight_inter_2_1_rdy),
      .weight_in_msg(weight_inter_2_1_msg),
      .act_in_val(act_inter_3_0_val),
      .act_in_rdy(act_inter_3_0_rdy),
      .act_in_msg(act_inter_3_0_msg),
      .accum_in_val(accum_inter_3_1_val),
      .accum_in_rdy(accum_inter_3_1_rdy),
      .accum_in_msg(accum_inter_3_1_msg),
      .weight_out_val(weight_inter_3_1_val),
      .weight_out_rdy(weight_inter_3_1_rdy),
      .weight_out_msg(weight_inter_3_1_msg),
      .act_out_val(act_inter_3_1_val),
      .act_out_rdy(act_inter_3_1_rdy),
      .act_out_msg(act_inter_3_1_msg),
      .accum_out_val(accum_inter_4_1_val),
      .accum_out_rdy(accum_inter_4_1_rdy),
      .accum_out_msg(accum_inter_4_1_msg)
    );
  SysPE SysPE_27 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_2_val),
      .weight_in_rdy(weight_inter_2_2_rdy),
      .weight_in_msg(weight_inter_2_2_msg),
      .act_in_val(act_inter_3_1_val),
      .act_in_rdy(act_inter_3_1_rdy),
      .act_in_msg(act_inter_3_1_msg),
      .accum_in_val(accum_inter_3_2_val),
      .accum_in_rdy(accum_inter_3_2_rdy),
      .accum_in_msg(accum_inter_3_2_msg),
      .weight_out_val(weight_inter_3_2_val),
      .weight_out_rdy(weight_inter_3_2_rdy),
      .weight_out_msg(weight_inter_3_2_msg),
      .act_out_val(act_inter_3_2_val),
      .act_out_rdy(act_inter_3_2_rdy),
      .act_out_msg(act_inter_3_2_msg),
      .accum_out_val(accum_inter_4_2_val),
      .accum_out_rdy(accum_inter_4_2_rdy),
      .accum_out_msg(accum_inter_4_2_msg)
    );
  SysPE SysPE_28 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_3_val),
      .weight_in_rdy(weight_inter_2_3_rdy),
      .weight_in_msg(weight_inter_2_3_msg),
      .act_in_val(act_inter_3_2_val),
      .act_in_rdy(act_inter_3_2_rdy),
      .act_in_msg(act_inter_3_2_msg),
      .accum_in_val(accum_inter_3_3_val),
      .accum_in_rdy(accum_inter_3_3_rdy),
      .accum_in_msg(accum_inter_3_3_msg),
      .weight_out_val(weight_inter_3_3_val),
      .weight_out_rdy(weight_inter_3_3_rdy),
      .weight_out_msg(weight_inter_3_3_msg),
      .act_out_val(act_inter_3_3_val),
      .act_out_rdy(act_inter_3_3_rdy),
      .act_out_msg(act_inter_3_3_msg),
      .accum_out_val(accum_inter_4_3_val),
      .accum_out_rdy(accum_inter_4_3_rdy),
      .accum_out_msg(accum_inter_4_3_msg)
    );
  SysPE SysPE_29 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_4_val),
      .weight_in_rdy(weight_inter_2_4_rdy),
      .weight_in_msg(weight_inter_2_4_msg),
      .act_in_val(act_inter_3_3_val),
      .act_in_rdy(act_inter_3_3_rdy),
      .act_in_msg(act_inter_3_3_msg),
      .accum_in_val(accum_inter_3_4_val),
      .accum_in_rdy(accum_inter_3_4_rdy),
      .accum_in_msg(accum_inter_3_4_msg),
      .weight_out_val(weight_inter_3_4_val),
      .weight_out_rdy(weight_inter_3_4_rdy),
      .weight_out_msg(weight_inter_3_4_msg),
      .act_out_val(act_inter_3_4_val),
      .act_out_rdy(act_inter_3_4_rdy),
      .act_out_msg(act_inter_3_4_msg),
      .accum_out_val(accum_inter_4_4_val),
      .accum_out_rdy(accum_inter_4_4_rdy),
      .accum_out_msg(accum_inter_4_4_msg)
    );
  SysPE SysPE_30 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_5_val),
      .weight_in_rdy(weight_inter_2_5_rdy),
      .weight_in_msg(weight_inter_2_5_msg),
      .act_in_val(act_inter_3_4_val),
      .act_in_rdy(act_inter_3_4_rdy),
      .act_in_msg(act_inter_3_4_msg),
      .accum_in_val(accum_inter_3_5_val),
      .accum_in_rdy(accum_inter_3_5_rdy),
      .accum_in_msg(accum_inter_3_5_msg),
      .weight_out_val(weight_inter_3_5_val),
      .weight_out_rdy(weight_inter_3_5_rdy),
      .weight_out_msg(weight_inter_3_5_msg),
      .act_out_val(act_inter_3_5_val),
      .act_out_rdy(act_inter_3_5_rdy),
      .act_out_msg(act_inter_3_5_msg),
      .accum_out_val(accum_inter_4_5_val),
      .accum_out_rdy(accum_inter_4_5_rdy),
      .accum_out_msg(accum_inter_4_5_msg)
    );
  SysPE SysPE_31 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_6_val),
      .weight_in_rdy(weight_inter_2_6_rdy),
      .weight_in_msg(weight_inter_2_6_msg),
      .act_in_val(act_inter_3_5_val),
      .act_in_rdy(act_inter_3_5_rdy),
      .act_in_msg(act_inter_3_5_msg),
      .accum_in_val(accum_inter_3_6_val),
      .accum_in_rdy(accum_inter_3_6_rdy),
      .accum_in_msg(accum_inter_3_6_msg),
      .weight_out_val(weight_inter_3_6_val),
      .weight_out_rdy(weight_inter_3_6_rdy),
      .weight_out_msg(weight_inter_3_6_msg),
      .act_out_val(act_inter_3_6_val),
      .act_out_rdy(act_inter_3_6_rdy),
      .act_out_msg(act_inter_3_6_msg),
      .accum_out_val(accum_inter_4_6_val),
      .accum_out_rdy(accum_inter_4_6_rdy),
      .accum_out_msg(accum_inter_4_6_msg)
    );
  SysPE SysPE_32 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_7_val),
      .weight_in_rdy(weight_inter_2_7_rdy),
      .weight_in_msg(weight_inter_2_7_msg),
      .act_in_val(act_inter_3_6_val),
      .act_in_rdy(act_inter_3_6_rdy),
      .act_in_msg(act_inter_3_6_msg),
      .accum_in_val(accum_inter_3_7_val),
      .accum_in_rdy(accum_inter_3_7_rdy),
      .accum_in_msg(accum_inter_3_7_msg),
      .weight_out_val(weight_inter_3_7_val),
      .weight_out_rdy(weight_inter_3_7_rdy),
      .weight_out_msg(weight_inter_3_7_msg),
      .act_out_val(act_inter_3_7_val),
      .act_out_rdy(act_inter_3_7_rdy),
      .act_out_msg(act_inter_3_7_msg),
      .accum_out_val(accum_inter_4_7_val),
      .accum_out_rdy(accum_inter_4_7_rdy),
      .accum_out_msg(accum_inter_4_7_msg)
    );
  SysPE SysPE_33 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_0_val),
      .weight_in_rdy(weight_inter_3_0_rdy),
      .weight_in_msg(weight_inter_3_0_msg),
      .act_in_val(act_in_vec_4_val),
      .act_in_rdy(act_in_vec_4_rdy),
      .act_in_msg(act_in_vec_4_msg),
      .accum_in_val(accum_inter_4_0_val),
      .accum_in_rdy(accum_inter_4_0_rdy),
      .accum_in_msg(accum_inter_4_0_msg),
      .weight_out_val(weight_inter_4_0_val),
      .weight_out_rdy(weight_inter_4_0_rdy),
      .weight_out_msg(weight_inter_4_0_msg),
      .act_out_val(act_inter_4_0_val),
      .act_out_rdy(act_inter_4_0_rdy),
      .act_out_msg(act_inter_4_0_msg),
      .accum_out_val(accum_inter_5_0_val),
      .accum_out_rdy(accum_inter_5_0_rdy),
      .accum_out_msg(accum_inter_5_0_msg)
    );
  SysPE SysPE_34 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_1_val),
      .weight_in_rdy(weight_inter_3_1_rdy),
      .weight_in_msg(weight_inter_3_1_msg),
      .act_in_val(act_inter_4_0_val),
      .act_in_rdy(act_inter_4_0_rdy),
      .act_in_msg(act_inter_4_0_msg),
      .accum_in_val(accum_inter_4_1_val),
      .accum_in_rdy(accum_inter_4_1_rdy),
      .accum_in_msg(accum_inter_4_1_msg),
      .weight_out_val(weight_inter_4_1_val),
      .weight_out_rdy(weight_inter_4_1_rdy),
      .weight_out_msg(weight_inter_4_1_msg),
      .act_out_val(act_inter_4_1_val),
      .act_out_rdy(act_inter_4_1_rdy),
      .act_out_msg(act_inter_4_1_msg),
      .accum_out_val(accum_inter_5_1_val),
      .accum_out_rdy(accum_inter_5_1_rdy),
      .accum_out_msg(accum_inter_5_1_msg)
    );
  SysPE SysPE_35 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_2_val),
      .weight_in_rdy(weight_inter_3_2_rdy),
      .weight_in_msg(weight_inter_3_2_msg),
      .act_in_val(act_inter_4_1_val),
      .act_in_rdy(act_inter_4_1_rdy),
      .act_in_msg(act_inter_4_1_msg),
      .accum_in_val(accum_inter_4_2_val),
      .accum_in_rdy(accum_inter_4_2_rdy),
      .accum_in_msg(accum_inter_4_2_msg),
      .weight_out_val(weight_inter_4_2_val),
      .weight_out_rdy(weight_inter_4_2_rdy),
      .weight_out_msg(weight_inter_4_2_msg),
      .act_out_val(act_inter_4_2_val),
      .act_out_rdy(act_inter_4_2_rdy),
      .act_out_msg(act_inter_4_2_msg),
      .accum_out_val(accum_inter_5_2_val),
      .accum_out_rdy(accum_inter_5_2_rdy),
      .accum_out_msg(accum_inter_5_2_msg)
    );
  SysPE SysPE_36 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_3_val),
      .weight_in_rdy(weight_inter_3_3_rdy),
      .weight_in_msg(weight_inter_3_3_msg),
      .act_in_val(act_inter_4_2_val),
      .act_in_rdy(act_inter_4_2_rdy),
      .act_in_msg(act_inter_4_2_msg),
      .accum_in_val(accum_inter_4_3_val),
      .accum_in_rdy(accum_inter_4_3_rdy),
      .accum_in_msg(accum_inter_4_3_msg),
      .weight_out_val(weight_inter_4_3_val),
      .weight_out_rdy(weight_inter_4_3_rdy),
      .weight_out_msg(weight_inter_4_3_msg),
      .act_out_val(act_inter_4_3_val),
      .act_out_rdy(act_inter_4_3_rdy),
      .act_out_msg(act_inter_4_3_msg),
      .accum_out_val(accum_inter_5_3_val),
      .accum_out_rdy(accum_inter_5_3_rdy),
      .accum_out_msg(accum_inter_5_3_msg)
    );
  SysPE SysPE_37 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_4_val),
      .weight_in_rdy(weight_inter_3_4_rdy),
      .weight_in_msg(weight_inter_3_4_msg),
      .act_in_val(act_inter_4_3_val),
      .act_in_rdy(act_inter_4_3_rdy),
      .act_in_msg(act_inter_4_3_msg),
      .accum_in_val(accum_inter_4_4_val),
      .accum_in_rdy(accum_inter_4_4_rdy),
      .accum_in_msg(accum_inter_4_4_msg),
      .weight_out_val(weight_inter_4_4_val),
      .weight_out_rdy(weight_inter_4_4_rdy),
      .weight_out_msg(weight_inter_4_4_msg),
      .act_out_val(act_inter_4_4_val),
      .act_out_rdy(act_inter_4_4_rdy),
      .act_out_msg(act_inter_4_4_msg),
      .accum_out_val(accum_inter_5_4_val),
      .accum_out_rdy(accum_inter_5_4_rdy),
      .accum_out_msg(accum_inter_5_4_msg)
    );
  SysPE SysPE_38 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_5_val),
      .weight_in_rdy(weight_inter_3_5_rdy),
      .weight_in_msg(weight_inter_3_5_msg),
      .act_in_val(act_inter_4_4_val),
      .act_in_rdy(act_inter_4_4_rdy),
      .act_in_msg(act_inter_4_4_msg),
      .accum_in_val(accum_inter_4_5_val),
      .accum_in_rdy(accum_inter_4_5_rdy),
      .accum_in_msg(accum_inter_4_5_msg),
      .weight_out_val(weight_inter_4_5_val),
      .weight_out_rdy(weight_inter_4_5_rdy),
      .weight_out_msg(weight_inter_4_5_msg),
      .act_out_val(act_inter_4_5_val),
      .act_out_rdy(act_inter_4_5_rdy),
      .act_out_msg(act_inter_4_5_msg),
      .accum_out_val(accum_inter_5_5_val),
      .accum_out_rdy(accum_inter_5_5_rdy),
      .accum_out_msg(accum_inter_5_5_msg)
    );
  SysPE SysPE_39 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_6_val),
      .weight_in_rdy(weight_inter_3_6_rdy),
      .weight_in_msg(weight_inter_3_6_msg),
      .act_in_val(act_inter_4_5_val),
      .act_in_rdy(act_inter_4_5_rdy),
      .act_in_msg(act_inter_4_5_msg),
      .accum_in_val(accum_inter_4_6_val),
      .accum_in_rdy(accum_inter_4_6_rdy),
      .accum_in_msg(accum_inter_4_6_msg),
      .weight_out_val(weight_inter_4_6_val),
      .weight_out_rdy(weight_inter_4_6_rdy),
      .weight_out_msg(weight_inter_4_6_msg),
      .act_out_val(act_inter_4_6_val),
      .act_out_rdy(act_inter_4_6_rdy),
      .act_out_msg(act_inter_4_6_msg),
      .accum_out_val(accum_inter_5_6_val),
      .accum_out_rdy(accum_inter_5_6_rdy),
      .accum_out_msg(accum_inter_5_6_msg)
    );
  SysPE SysPE_40 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_7_val),
      .weight_in_rdy(weight_inter_3_7_rdy),
      .weight_in_msg(weight_inter_3_7_msg),
      .act_in_val(act_inter_4_6_val),
      .act_in_rdy(act_inter_4_6_rdy),
      .act_in_msg(act_inter_4_6_msg),
      .accum_in_val(accum_inter_4_7_val),
      .accum_in_rdy(accum_inter_4_7_rdy),
      .accum_in_msg(accum_inter_4_7_msg),
      .weight_out_val(weight_inter_4_7_val),
      .weight_out_rdy(weight_inter_4_7_rdy),
      .weight_out_msg(weight_inter_4_7_msg),
      .act_out_val(act_inter_4_7_val),
      .act_out_rdy(act_inter_4_7_rdy),
      .act_out_msg(act_inter_4_7_msg),
      .accum_out_val(accum_inter_5_7_val),
      .accum_out_rdy(accum_inter_5_7_rdy),
      .accum_out_msg(accum_inter_5_7_msg)
    );
  SysPE SysPE_41 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_0_val),
      .weight_in_rdy(weight_inter_4_0_rdy),
      .weight_in_msg(weight_inter_4_0_msg),
      .act_in_val(act_in_vec_5_val),
      .act_in_rdy(act_in_vec_5_rdy),
      .act_in_msg(act_in_vec_5_msg),
      .accum_in_val(accum_inter_5_0_val),
      .accum_in_rdy(accum_inter_5_0_rdy),
      .accum_in_msg(accum_inter_5_0_msg),
      .weight_out_val(weight_inter_5_0_val),
      .weight_out_rdy(weight_inter_5_0_rdy),
      .weight_out_msg(weight_inter_5_0_msg),
      .act_out_val(act_inter_5_0_val),
      .act_out_rdy(act_inter_5_0_rdy),
      .act_out_msg(act_inter_5_0_msg),
      .accum_out_val(accum_inter_6_0_val),
      .accum_out_rdy(accum_inter_6_0_rdy),
      .accum_out_msg(accum_inter_6_0_msg)
    );
  SysPE SysPE_42 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_1_val),
      .weight_in_rdy(weight_inter_4_1_rdy),
      .weight_in_msg(weight_inter_4_1_msg),
      .act_in_val(act_inter_5_0_val),
      .act_in_rdy(act_inter_5_0_rdy),
      .act_in_msg(act_inter_5_0_msg),
      .accum_in_val(accum_inter_5_1_val),
      .accum_in_rdy(accum_inter_5_1_rdy),
      .accum_in_msg(accum_inter_5_1_msg),
      .weight_out_val(weight_inter_5_1_val),
      .weight_out_rdy(weight_inter_5_1_rdy),
      .weight_out_msg(weight_inter_5_1_msg),
      .act_out_val(act_inter_5_1_val),
      .act_out_rdy(act_inter_5_1_rdy),
      .act_out_msg(act_inter_5_1_msg),
      .accum_out_val(accum_inter_6_1_val),
      .accum_out_rdy(accum_inter_6_1_rdy),
      .accum_out_msg(accum_inter_6_1_msg)
    );
  SysPE SysPE_43 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_2_val),
      .weight_in_rdy(weight_inter_4_2_rdy),
      .weight_in_msg(weight_inter_4_2_msg),
      .act_in_val(act_inter_5_1_val),
      .act_in_rdy(act_inter_5_1_rdy),
      .act_in_msg(act_inter_5_1_msg),
      .accum_in_val(accum_inter_5_2_val),
      .accum_in_rdy(accum_inter_5_2_rdy),
      .accum_in_msg(accum_inter_5_2_msg),
      .weight_out_val(weight_inter_5_2_val),
      .weight_out_rdy(weight_inter_5_2_rdy),
      .weight_out_msg(weight_inter_5_2_msg),
      .act_out_val(act_inter_5_2_val),
      .act_out_rdy(act_inter_5_2_rdy),
      .act_out_msg(act_inter_5_2_msg),
      .accum_out_val(accum_inter_6_2_val),
      .accum_out_rdy(accum_inter_6_2_rdy),
      .accum_out_msg(accum_inter_6_2_msg)
    );
  SysPE SysPE_44 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_3_val),
      .weight_in_rdy(weight_inter_4_3_rdy),
      .weight_in_msg(weight_inter_4_3_msg),
      .act_in_val(act_inter_5_2_val),
      .act_in_rdy(act_inter_5_2_rdy),
      .act_in_msg(act_inter_5_2_msg),
      .accum_in_val(accum_inter_5_3_val),
      .accum_in_rdy(accum_inter_5_3_rdy),
      .accum_in_msg(accum_inter_5_3_msg),
      .weight_out_val(weight_inter_5_3_val),
      .weight_out_rdy(weight_inter_5_3_rdy),
      .weight_out_msg(weight_inter_5_3_msg),
      .act_out_val(act_inter_5_3_val),
      .act_out_rdy(act_inter_5_3_rdy),
      .act_out_msg(act_inter_5_3_msg),
      .accum_out_val(accum_inter_6_3_val),
      .accum_out_rdy(accum_inter_6_3_rdy),
      .accum_out_msg(accum_inter_6_3_msg)
    );
  SysPE SysPE_45 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_4_val),
      .weight_in_rdy(weight_inter_4_4_rdy),
      .weight_in_msg(weight_inter_4_4_msg),
      .act_in_val(act_inter_5_3_val),
      .act_in_rdy(act_inter_5_3_rdy),
      .act_in_msg(act_inter_5_3_msg),
      .accum_in_val(accum_inter_5_4_val),
      .accum_in_rdy(accum_inter_5_4_rdy),
      .accum_in_msg(accum_inter_5_4_msg),
      .weight_out_val(weight_inter_5_4_val),
      .weight_out_rdy(weight_inter_5_4_rdy),
      .weight_out_msg(weight_inter_5_4_msg),
      .act_out_val(act_inter_5_4_val),
      .act_out_rdy(act_inter_5_4_rdy),
      .act_out_msg(act_inter_5_4_msg),
      .accum_out_val(accum_inter_6_4_val),
      .accum_out_rdy(accum_inter_6_4_rdy),
      .accum_out_msg(accum_inter_6_4_msg)
    );
  SysPE SysPE_46 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_5_val),
      .weight_in_rdy(weight_inter_4_5_rdy),
      .weight_in_msg(weight_inter_4_5_msg),
      .act_in_val(act_inter_5_4_val),
      .act_in_rdy(act_inter_5_4_rdy),
      .act_in_msg(act_inter_5_4_msg),
      .accum_in_val(accum_inter_5_5_val),
      .accum_in_rdy(accum_inter_5_5_rdy),
      .accum_in_msg(accum_inter_5_5_msg),
      .weight_out_val(weight_inter_5_5_val),
      .weight_out_rdy(weight_inter_5_5_rdy),
      .weight_out_msg(weight_inter_5_5_msg),
      .act_out_val(act_inter_5_5_val),
      .act_out_rdy(act_inter_5_5_rdy),
      .act_out_msg(act_inter_5_5_msg),
      .accum_out_val(accum_inter_6_5_val),
      .accum_out_rdy(accum_inter_6_5_rdy),
      .accum_out_msg(accum_inter_6_5_msg)
    );
  SysPE SysPE_47 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_6_val),
      .weight_in_rdy(weight_inter_4_6_rdy),
      .weight_in_msg(weight_inter_4_6_msg),
      .act_in_val(act_inter_5_5_val),
      .act_in_rdy(act_inter_5_5_rdy),
      .act_in_msg(act_inter_5_5_msg),
      .accum_in_val(accum_inter_5_6_val),
      .accum_in_rdy(accum_inter_5_6_rdy),
      .accum_in_msg(accum_inter_5_6_msg),
      .weight_out_val(weight_inter_5_6_val),
      .weight_out_rdy(weight_inter_5_6_rdy),
      .weight_out_msg(weight_inter_5_6_msg),
      .act_out_val(act_inter_5_6_val),
      .act_out_rdy(act_inter_5_6_rdy),
      .act_out_msg(act_inter_5_6_msg),
      .accum_out_val(accum_inter_6_6_val),
      .accum_out_rdy(accum_inter_6_6_rdy),
      .accum_out_msg(accum_inter_6_6_msg)
    );
  SysPE SysPE_48 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_7_val),
      .weight_in_rdy(weight_inter_4_7_rdy),
      .weight_in_msg(weight_inter_4_7_msg),
      .act_in_val(act_inter_5_6_val),
      .act_in_rdy(act_inter_5_6_rdy),
      .act_in_msg(act_inter_5_6_msg),
      .accum_in_val(accum_inter_5_7_val),
      .accum_in_rdy(accum_inter_5_7_rdy),
      .accum_in_msg(accum_inter_5_7_msg),
      .weight_out_val(weight_inter_5_7_val),
      .weight_out_rdy(weight_inter_5_7_rdy),
      .weight_out_msg(weight_inter_5_7_msg),
      .act_out_val(act_inter_5_7_val),
      .act_out_rdy(act_inter_5_7_rdy),
      .act_out_msg(act_inter_5_7_msg),
      .accum_out_val(accum_inter_6_7_val),
      .accum_out_rdy(accum_inter_6_7_rdy),
      .accum_out_msg(accum_inter_6_7_msg)
    );
  SysPE SysPE_49 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_0_val),
      .weight_in_rdy(weight_inter_5_0_rdy),
      .weight_in_msg(weight_inter_5_0_msg),
      .act_in_val(act_in_vec_6_val),
      .act_in_rdy(act_in_vec_6_rdy),
      .act_in_msg(act_in_vec_6_msg),
      .accum_in_val(accum_inter_6_0_val),
      .accum_in_rdy(accum_inter_6_0_rdy),
      .accum_in_msg(accum_inter_6_0_msg),
      .weight_out_val(weight_inter_6_0_val),
      .weight_out_rdy(weight_inter_6_0_rdy),
      .weight_out_msg(weight_inter_6_0_msg),
      .act_out_val(act_inter_6_0_val),
      .act_out_rdy(act_inter_6_0_rdy),
      .act_out_msg(act_inter_6_0_msg),
      .accum_out_val(accum_inter_7_0_val),
      .accum_out_rdy(accum_inter_7_0_rdy),
      .accum_out_msg(accum_inter_7_0_msg)
    );
  SysPE SysPE_50 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_1_val),
      .weight_in_rdy(weight_inter_5_1_rdy),
      .weight_in_msg(weight_inter_5_1_msg),
      .act_in_val(act_inter_6_0_val),
      .act_in_rdy(act_inter_6_0_rdy),
      .act_in_msg(act_inter_6_0_msg),
      .accum_in_val(accum_inter_6_1_val),
      .accum_in_rdy(accum_inter_6_1_rdy),
      .accum_in_msg(accum_inter_6_1_msg),
      .weight_out_val(weight_inter_6_1_val),
      .weight_out_rdy(weight_inter_6_1_rdy),
      .weight_out_msg(weight_inter_6_1_msg),
      .act_out_val(act_inter_6_1_val),
      .act_out_rdy(act_inter_6_1_rdy),
      .act_out_msg(act_inter_6_1_msg),
      .accum_out_val(accum_inter_7_1_val),
      .accum_out_rdy(accum_inter_7_1_rdy),
      .accum_out_msg(accum_inter_7_1_msg)
    );
  SysPE SysPE_51 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_2_val),
      .weight_in_rdy(weight_inter_5_2_rdy),
      .weight_in_msg(weight_inter_5_2_msg),
      .act_in_val(act_inter_6_1_val),
      .act_in_rdy(act_inter_6_1_rdy),
      .act_in_msg(act_inter_6_1_msg),
      .accum_in_val(accum_inter_6_2_val),
      .accum_in_rdy(accum_inter_6_2_rdy),
      .accum_in_msg(accum_inter_6_2_msg),
      .weight_out_val(weight_inter_6_2_val),
      .weight_out_rdy(weight_inter_6_2_rdy),
      .weight_out_msg(weight_inter_6_2_msg),
      .act_out_val(act_inter_6_2_val),
      .act_out_rdy(act_inter_6_2_rdy),
      .act_out_msg(act_inter_6_2_msg),
      .accum_out_val(accum_inter_7_2_val),
      .accum_out_rdy(accum_inter_7_2_rdy),
      .accum_out_msg(accum_inter_7_2_msg)
    );
  SysPE SysPE_52 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_3_val),
      .weight_in_rdy(weight_inter_5_3_rdy),
      .weight_in_msg(weight_inter_5_3_msg),
      .act_in_val(act_inter_6_2_val),
      .act_in_rdy(act_inter_6_2_rdy),
      .act_in_msg(act_inter_6_2_msg),
      .accum_in_val(accum_inter_6_3_val),
      .accum_in_rdy(accum_inter_6_3_rdy),
      .accum_in_msg(accum_inter_6_3_msg),
      .weight_out_val(weight_inter_6_3_val),
      .weight_out_rdy(weight_inter_6_3_rdy),
      .weight_out_msg(weight_inter_6_3_msg),
      .act_out_val(act_inter_6_3_val),
      .act_out_rdy(act_inter_6_3_rdy),
      .act_out_msg(act_inter_6_3_msg),
      .accum_out_val(accum_inter_7_3_val),
      .accum_out_rdy(accum_inter_7_3_rdy),
      .accum_out_msg(accum_inter_7_3_msg)
    );
  SysPE SysPE_53 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_4_val),
      .weight_in_rdy(weight_inter_5_4_rdy),
      .weight_in_msg(weight_inter_5_4_msg),
      .act_in_val(act_inter_6_3_val),
      .act_in_rdy(act_inter_6_3_rdy),
      .act_in_msg(act_inter_6_3_msg),
      .accum_in_val(accum_inter_6_4_val),
      .accum_in_rdy(accum_inter_6_4_rdy),
      .accum_in_msg(accum_inter_6_4_msg),
      .weight_out_val(weight_inter_6_4_val),
      .weight_out_rdy(weight_inter_6_4_rdy),
      .weight_out_msg(weight_inter_6_4_msg),
      .act_out_val(act_inter_6_4_val),
      .act_out_rdy(act_inter_6_4_rdy),
      .act_out_msg(act_inter_6_4_msg),
      .accum_out_val(accum_inter_7_4_val),
      .accum_out_rdy(accum_inter_7_4_rdy),
      .accum_out_msg(accum_inter_7_4_msg)
    );
  SysPE SysPE_54 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_5_val),
      .weight_in_rdy(weight_inter_5_5_rdy),
      .weight_in_msg(weight_inter_5_5_msg),
      .act_in_val(act_inter_6_4_val),
      .act_in_rdy(act_inter_6_4_rdy),
      .act_in_msg(act_inter_6_4_msg),
      .accum_in_val(accum_inter_6_5_val),
      .accum_in_rdy(accum_inter_6_5_rdy),
      .accum_in_msg(accum_inter_6_5_msg),
      .weight_out_val(weight_inter_6_5_val),
      .weight_out_rdy(weight_inter_6_5_rdy),
      .weight_out_msg(weight_inter_6_5_msg),
      .act_out_val(act_inter_6_5_val),
      .act_out_rdy(act_inter_6_5_rdy),
      .act_out_msg(act_inter_6_5_msg),
      .accum_out_val(accum_inter_7_5_val),
      .accum_out_rdy(accum_inter_7_5_rdy),
      .accum_out_msg(accum_inter_7_5_msg)
    );
  SysPE SysPE_55 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_6_val),
      .weight_in_rdy(weight_inter_5_6_rdy),
      .weight_in_msg(weight_inter_5_6_msg),
      .act_in_val(act_inter_6_5_val),
      .act_in_rdy(act_inter_6_5_rdy),
      .act_in_msg(act_inter_6_5_msg),
      .accum_in_val(accum_inter_6_6_val),
      .accum_in_rdy(accum_inter_6_6_rdy),
      .accum_in_msg(accum_inter_6_6_msg),
      .weight_out_val(weight_inter_6_6_val),
      .weight_out_rdy(weight_inter_6_6_rdy),
      .weight_out_msg(weight_inter_6_6_msg),
      .act_out_val(act_inter_6_6_val),
      .act_out_rdy(act_inter_6_6_rdy),
      .act_out_msg(act_inter_6_6_msg),
      .accum_out_val(accum_inter_7_6_val),
      .accum_out_rdy(accum_inter_7_6_rdy),
      .accum_out_msg(accum_inter_7_6_msg)
    );
  SysPE SysPE_56 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_7_val),
      .weight_in_rdy(weight_inter_5_7_rdy),
      .weight_in_msg(weight_inter_5_7_msg),
      .act_in_val(act_inter_6_6_val),
      .act_in_rdy(act_inter_6_6_rdy),
      .act_in_msg(act_inter_6_6_msg),
      .accum_in_val(accum_inter_6_7_val),
      .accum_in_rdy(accum_inter_6_7_rdy),
      .accum_in_msg(accum_inter_6_7_msg),
      .weight_out_val(weight_inter_6_7_val),
      .weight_out_rdy(weight_inter_6_7_rdy),
      .weight_out_msg(weight_inter_6_7_msg),
      .act_out_val(act_inter_6_7_val),
      .act_out_rdy(act_inter_6_7_rdy),
      .act_out_msg(act_inter_6_7_msg),
      .accum_out_val(accum_inter_7_7_val),
      .accum_out_rdy(accum_inter_7_7_rdy),
      .accum_out_msg(accum_inter_7_7_msg)
    );
  SysPE SysPE_57 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_0_val),
      .weight_in_rdy(weight_inter_6_0_rdy),
      .weight_in_msg(weight_inter_6_0_msg),
      .act_in_val(act_in_vec_7_val),
      .act_in_rdy(act_in_vec_7_rdy),
      .act_in_msg(act_in_vec_7_msg),
      .accum_in_val(accum_inter_7_0_val),
      .accum_in_rdy(accum_inter_7_0_rdy),
      .accum_in_msg(accum_inter_7_0_msg),
      .weight_out_val(weight_inter_7_0_val),
      .weight_out_rdy(weight_inter_7_0_rdy),
      .weight_out_msg(weight_inter_7_0_msg),
      .act_out_val(act_inter_7_0_val),
      .act_out_rdy(act_inter_7_0_rdy),
      .act_out_msg(act_inter_7_0_msg),
      .accum_out_val(accum_out_vec_0_val),
      .accum_out_rdy(accum_out_vec_0_rdy),
      .accum_out_msg(accum_out_vec_0_msg)
    );
  SysPE SysPE_58 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_1_val),
      .weight_in_rdy(weight_inter_6_1_rdy),
      .weight_in_msg(weight_inter_6_1_msg),
      .act_in_val(act_inter_7_0_val),
      .act_in_rdy(act_inter_7_0_rdy),
      .act_in_msg(act_inter_7_0_msg),
      .accum_in_val(accum_inter_7_1_val),
      .accum_in_rdy(accum_inter_7_1_rdy),
      .accum_in_msg(accum_inter_7_1_msg),
      .weight_out_val(weight_inter_7_1_val),
      .weight_out_rdy(weight_inter_7_1_rdy),
      .weight_out_msg(weight_inter_7_1_msg),
      .act_out_val(act_inter_7_1_val),
      .act_out_rdy(act_inter_7_1_rdy),
      .act_out_msg(act_inter_7_1_msg),
      .accum_out_val(accum_out_vec_1_val),
      .accum_out_rdy(accum_out_vec_1_rdy),
      .accum_out_msg(accum_out_vec_1_msg)
    );
  SysPE SysPE_59 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_2_val),
      .weight_in_rdy(weight_inter_6_2_rdy),
      .weight_in_msg(weight_inter_6_2_msg),
      .act_in_val(act_inter_7_1_val),
      .act_in_rdy(act_inter_7_1_rdy),
      .act_in_msg(act_inter_7_1_msg),
      .accum_in_val(accum_inter_7_2_val),
      .accum_in_rdy(accum_inter_7_2_rdy),
      .accum_in_msg(accum_inter_7_2_msg),
      .weight_out_val(weight_inter_7_2_val),
      .weight_out_rdy(weight_inter_7_2_rdy),
      .weight_out_msg(weight_inter_7_2_msg),
      .act_out_val(act_inter_7_2_val),
      .act_out_rdy(act_inter_7_2_rdy),
      .act_out_msg(act_inter_7_2_msg),
      .accum_out_val(accum_out_vec_2_val),
      .accum_out_rdy(accum_out_vec_2_rdy),
      .accum_out_msg(accum_out_vec_2_msg)
    );
  SysPE SysPE_60 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_3_val),
      .weight_in_rdy(weight_inter_6_3_rdy),
      .weight_in_msg(weight_inter_6_3_msg),
      .act_in_val(act_inter_7_2_val),
      .act_in_rdy(act_inter_7_2_rdy),
      .act_in_msg(act_inter_7_2_msg),
      .accum_in_val(accum_inter_7_3_val),
      .accum_in_rdy(accum_inter_7_3_rdy),
      .accum_in_msg(accum_inter_7_3_msg),
      .weight_out_val(weight_inter_7_3_val),
      .weight_out_rdy(weight_inter_7_3_rdy),
      .weight_out_msg(weight_inter_7_3_msg),
      .act_out_val(act_inter_7_3_val),
      .act_out_rdy(act_inter_7_3_rdy),
      .act_out_msg(act_inter_7_3_msg),
      .accum_out_val(accum_out_vec_3_val),
      .accum_out_rdy(accum_out_vec_3_rdy),
      .accum_out_msg(accum_out_vec_3_msg)
    );
  SysPE SysPE_61 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_4_val),
      .weight_in_rdy(weight_inter_6_4_rdy),
      .weight_in_msg(weight_inter_6_4_msg),
      .act_in_val(act_inter_7_3_val),
      .act_in_rdy(act_inter_7_3_rdy),
      .act_in_msg(act_inter_7_3_msg),
      .accum_in_val(accum_inter_7_4_val),
      .accum_in_rdy(accum_inter_7_4_rdy),
      .accum_in_msg(accum_inter_7_4_msg),
      .weight_out_val(weight_inter_7_4_val),
      .weight_out_rdy(weight_inter_7_4_rdy),
      .weight_out_msg(weight_inter_7_4_msg),
      .act_out_val(act_inter_7_4_val),
      .act_out_rdy(act_inter_7_4_rdy),
      .act_out_msg(act_inter_7_4_msg),
      .accum_out_val(accum_out_vec_4_val),
      .accum_out_rdy(accum_out_vec_4_rdy),
      .accum_out_msg(accum_out_vec_4_msg)
    );
  SysPE SysPE_62 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_5_val),
      .weight_in_rdy(weight_inter_6_5_rdy),
      .weight_in_msg(weight_inter_6_5_msg),
      .act_in_val(act_inter_7_4_val),
      .act_in_rdy(act_inter_7_4_rdy),
      .act_in_msg(act_inter_7_4_msg),
      .accum_in_val(accum_inter_7_5_val),
      .accum_in_rdy(accum_inter_7_5_rdy),
      .accum_in_msg(accum_inter_7_5_msg),
      .weight_out_val(weight_inter_7_5_val),
      .weight_out_rdy(weight_inter_7_5_rdy),
      .weight_out_msg(weight_inter_7_5_msg),
      .act_out_val(act_inter_7_5_val),
      .act_out_rdy(act_inter_7_5_rdy),
      .act_out_msg(act_inter_7_5_msg),
      .accum_out_val(accum_out_vec_5_val),
      .accum_out_rdy(accum_out_vec_5_rdy),
      .accum_out_msg(accum_out_vec_5_msg)
    );
  SysPE SysPE_63 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_6_val),
      .weight_in_rdy(weight_inter_6_6_rdy),
      .weight_in_msg(weight_inter_6_6_msg),
      .act_in_val(act_inter_7_5_val),
      .act_in_rdy(act_inter_7_5_rdy),
      .act_in_msg(act_inter_7_5_msg),
      .accum_in_val(accum_inter_7_6_val),
      .accum_in_rdy(accum_inter_7_6_rdy),
      .accum_in_msg(accum_inter_7_6_msg),
      .weight_out_val(weight_inter_7_6_val),
      .weight_out_rdy(weight_inter_7_6_rdy),
      .weight_out_msg(weight_inter_7_6_msg),
      .act_out_val(act_inter_7_6_val),
      .act_out_rdy(act_inter_7_6_rdy),
      .act_out_msg(act_inter_7_6_msg),
      .accum_out_val(accum_out_vec_6_val),
      .accum_out_rdy(accum_out_vec_6_rdy),
      .accum_out_msg(accum_out_vec_6_msg)
    );
  SysPE SysPE_64 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_7_val),
      .weight_in_rdy(weight_inter_6_7_rdy),
      .weight_in_msg(weight_inter_6_7_msg),
      .act_in_val(act_inter_7_6_val),
      .act_in_rdy(act_inter_7_6_rdy),
      .act_in_msg(act_inter_7_6_msg),
      .accum_in_val(accum_inter_7_7_val),
      .accum_in_rdy(accum_inter_7_7_rdy),
      .accum_in_msg(accum_inter_7_7_msg),
      .weight_out_val(weight_inter_7_7_val),
      .weight_out_rdy(weight_inter_7_7_rdy),
      .weight_out_msg(weight_inter_7_7_msg),
      .act_out_val(act_inter_7_7_val),
      .act_out_rdy(act_inter_7_7_rdy),
      .act_out_msg(act_inter_7_7_msg),
      .accum_out_val(accum_out_vec_7_val),
      .accum_out_rdy(accum_out_vec_7_rdy),
      .accum_out_msg(accum_out_vec_7_msg)
    );
  SysArray_WeightOutRun SysArray_WeightOutRun_inst (
      .clk(clk),
      .rst(rst),
      .weight_inter_7_0_val(weight_inter_7_0_val),
      .weight_inter_7_1_val(weight_inter_7_1_val),
      .weight_inter_7_2_val(weight_inter_7_2_val),
      .weight_inter_7_3_val(weight_inter_7_3_val),
      .weight_inter_7_4_val(weight_inter_7_4_val),
      .weight_inter_7_5_val(weight_inter_7_5_val),
      .weight_inter_7_6_val(weight_inter_7_6_val),
      .weight_inter_7_7_val(weight_inter_7_7_val),
      .weight_inter_7_0_rdy(weight_inter_7_0_rdy),
      .weight_inter_7_1_rdy(weight_inter_7_1_rdy),
      .weight_inter_7_2_rdy(weight_inter_7_2_rdy),
      .weight_inter_7_3_rdy(weight_inter_7_3_rdy),
      .weight_inter_7_4_rdy(weight_inter_7_4_rdy),
      .weight_inter_7_5_rdy(weight_inter_7_5_rdy),
      .weight_inter_7_6_rdy(weight_inter_7_6_rdy),
      .weight_inter_7_7_rdy(weight_inter_7_7_rdy),
      .weight_inter_7_0_msg(weight_inter_7_0_msg),
      .weight_inter_7_1_msg(weight_inter_7_1_msg),
      .weight_inter_7_2_msg(weight_inter_7_2_msg),
      .weight_inter_7_3_msg(weight_inter_7_3_msg),
      .weight_inter_7_4_msg(weight_inter_7_4_msg),
      .weight_inter_7_5_msg(weight_inter_7_5_msg),
      .weight_inter_7_6_msg(weight_inter_7_6_msg),
      .weight_inter_7_7_msg(weight_inter_7_7_msg)
    );
  SysArray_ActOutRun SysArray_ActOutRun_inst (
      .clk(clk),
      .rst(rst),
      .act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_pff(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  SysArray_AccumInRun SysArray_AccumInRun_inst (
      .clk(clk),
      .rst(rst),
      .accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_pff(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
endmodule



