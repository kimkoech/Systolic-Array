
//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ../td_ccore_solutions/Connections__InBlocking_SysPE__InputType_Connections__SYN_--_3d75a24542f9bd72f21738470c667f036340_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Thu Apr 16 13:53:00 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  mgc_out_dreg_v2 #(.rscid(32'sd1),
  .width(32'sd8)) data_rsci (
      .d(nl_data_rsci_d[7:0]),
      .z(data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd22),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, do_wait_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  input do_wait_rsc_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__OutBlocking_SysPE__InputType_Connections__SYN--_7961c91e828f28e6b31ea17763393cd662ff_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Thu Apr 16 13:52:59 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB_core
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB_core (
  this_val, this_rdy, this_msg, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [7:0] this_msg;
  reg [7:0] this_msg;
  input [7:0] m_rsc_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [7:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire or_dcpl;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd8)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_rdy),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd21),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign or_dcpl = ccs_ccore_start_rsci_idat | asn_itm_1;
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 8'b00000000;
      this_val <= 1'b0;
    end
    else if ( or_dcpl ) begin
      this_msg <= MUX_v_8_2_2(8'b00000000, m_rsci_idat, ccs_ccore_start_rsci_idat);
      this_val <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end

  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB (
  this_val, this_rdy, this_msg, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [7:0] this_msg;
  input [7:0] m_rsc_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB_core Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__InBlocking_SysPE__AccumType_Connections__SYN_--_fcc000cdee2bdbaf1af8321dad3e708762fd_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Thu Apr 16 13:52:57 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [31:0] this_msg;
  output [31:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  mgc_out_dreg_v2 #(.rscid(32'sd7),
  .width(32'sd32)) data_rsci (
      .d(nl_data_rsci_d[31:0]),
      .z(data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd9),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd20),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, do_wait_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [31:0] this_msg;
  output [31:0] data_rsc_z;
  input do_wait_rsc_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ../td_ccore_solutions/Connections__OutBlocking_SysPE__InputType_Connections__SYN--_027f1954845d044556c8243937c776375bcb_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Thu Apr 16 13:52:55 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [7:0] this_msg;
  reg [7:0] this_msg;
  input [7:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [7:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd10),
  .width(32'sd8)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd19),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd24)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 8'b00000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_msg <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [7:0] this_msg;
  input [7:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__OutBlocking_SysPE__AccumType_Connections__SYN--_2c1d8b870a5e6780c1a757ef891031fc5be9_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Thu Apr 16 13:52:53 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [31:0] this_msg;
  reg [31:0] this_msg;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [31:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd11),
  .width(32'sd32)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd18),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd23)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_msg <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [31:0] this_msg;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 21:42:14 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_PERun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysPE_PERun_PERun_fsm (
  clk, rst, PERun_wen, fsm_output
);
  input clk;
  input rst;
  input PERun_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysPE_PERun_PERun_fsm_1
  parameter
    PERun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysPE_PERun_PERun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // PERun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PERun_rlp_C_0;
    end
    else if ( PERun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_staller
// ------------------------------------------------------------------


module SysPE_PERun_staller (
  clk, rst, PERun_wen, PERun_wten, act_out_Push_mioi_wen_comp, accum_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PERun_wen;
  output PERun_wten;
  input act_out_Push_mioi_wen_comp;
  input accum_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PERun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PERun_wen = act_out_Push_mioi_wen_comp & accum_out_Push_mioi_wen_comp;
  assign PERun_wten = PERun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PERun_wten_reg <= 1'b0;
    end
    else begin
      PERun_wten_reg <= ~ PERun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp (
  clk, rst, accum_out_Push_mioi_oswt, accum_out_Push_mioi_wen_comp, accum_out_Push_mioi_biwt,
      accum_out_Push_mioi_bdwt, accum_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_wen_comp;
  input accum_out_Push_mioi_biwt;
  input accum_out_Push_mioi_bdwt;
  output accum_out_Push_mioi_bcwt;
  reg accum_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign accum_out_Push_mioi_wen_comp = (~ accum_out_Push_mioi_oswt) | accum_out_Push_mioi_biwt
      | accum_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      accum_out_Push_mioi_bcwt <= ~((~(accum_out_Push_mioi_bcwt | accum_out_Push_mioi_biwt))
          | accum_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl (
  PERun_wen, accum_out_Push_mioi_oswt, accum_out_Push_mioi_biwt, accum_out_Push_mioi_bdwt,
      accum_out_Push_mioi_bcwt, accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct,
      accum_out_Push_mioi_ccs_ccore_done_sync_vld, accum_out_Push_mioi_oswt_pff
);
  input PERun_wen;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_biwt;
  output accum_out_Push_mioi_bdwt;
  input accum_out_Push_mioi_bcwt;
  output accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input accum_out_Push_mioi_ccs_ccore_done_sync_vld;
  input accum_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accum_out_Push_mioi_bdwt = accum_out_Push_mioi_oswt & PERun_wen;
  assign accum_out_Push_mioi_biwt = accum_out_Push_mioi_oswt & (~ accum_out_Push_mioi_bcwt)
      & accum_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct = accum_out_Push_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp (
  clk, rst, act_out_Push_mioi_oswt, act_out_Push_mioi_wen_comp, act_out_Push_mioi_biwt,
      act_out_Push_mioi_bdwt, act_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_wen_comp;
  input act_out_Push_mioi_biwt;
  input act_out_Push_mioi_bdwt;
  output act_out_Push_mioi_bcwt;
  reg act_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_out_Push_mioi_wen_comp = (~ act_out_Push_mioi_oswt) | act_out_Push_mioi_biwt
      | act_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_out_Push_mioi_bcwt <= ~((~(act_out_Push_mioi_bcwt | act_out_Push_mioi_biwt))
          | act_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl (
  PERun_wen, act_out_Push_mioi_oswt, act_out_Push_mioi_biwt, act_out_Push_mioi_bdwt,
      act_out_Push_mioi_bcwt, act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct,
      act_out_Push_mioi_ccs_ccore_done_sync_vld, act_out_Push_mioi_oswt_pff
);
  input PERun_wen;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_biwt;
  output act_out_Push_mioi_bdwt;
  input act_out_Push_mioi_bcwt;
  output act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input act_out_Push_mioi_ccs_ccore_done_sync_vld;
  input act_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_out_Push_mioi_bdwt = act_out_Push_mioi_oswt & PERun_wen;
  assign act_out_Push_mioi_biwt = act_out_Push_mioi_oswt & (~ act_out_Push_mioi_bcwt)
      & act_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct = act_out_Push_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp (
  clk, rst, accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_in_PopNB_mioi_return_rsc_z_mxwt,
      accum_in_PopNB_mioi_data_rsc_z, accum_in_PopNB_mioi_biwt, accum_in_PopNB_mioi_bdwt,
      accum_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  output accum_in_PopNB_mioi_return_rsc_z_mxwt;
  input [31:0] accum_in_PopNB_mioi_data_rsc_z;
  input accum_in_PopNB_mioi_biwt;
  input accum_in_PopNB_mioi_bdwt;
  input accum_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg accum_in_PopNB_mioi_bcwt;
  reg [31:0] accum_in_PopNB_mioi_data_rsc_z_bfwt;
  reg accum_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accum_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_32_2_2(accum_in_PopNB_mioi_data_rsc_z,
      accum_in_PopNB_mioi_data_rsc_z_bfwt, accum_in_PopNB_mioi_bcwt);
  assign accum_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(accum_in_PopNB_mioi_return_rsc_z,
      accum_in_PopNB_mioi_return_rsc_z_bfwt, accum_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_in_PopNB_mioi_bcwt <= 1'b0;
      accum_in_PopNB_mioi_data_rsc_z_bfwt <= 32'b00000000000000000000000000000000;
      accum_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      accum_in_PopNB_mioi_bcwt <= ~((~(accum_in_PopNB_mioi_bcwt | accum_in_PopNB_mioi_biwt))
          | accum_in_PopNB_mioi_bdwt);
      accum_in_PopNB_mioi_data_rsc_z_bfwt <= accum_in_PopNB_mioi_data_rsc_z_mxwt;
      accum_in_PopNB_mioi_return_rsc_z_bfwt <= accum_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl (
  PERun_wen, PERun_wten, accum_in_PopNB_mioi_oswt, accum_in_PopNB_mioi_biwt, accum_in_PopNB_mioi_bdwt,
      accum_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff, accum_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input PERun_wten;
  input accum_in_PopNB_mioi_oswt;
  output accum_in_PopNB_mioi_biwt;
  output accum_in_PopNB_mioi_bdwt;
  output accum_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff;
  input accum_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accum_in_PopNB_mioi_bdwt = accum_in_PopNB_mioi_oswt & PERun_wen;
  assign accum_in_PopNB_mioi_biwt = (~ PERun_wten) & accum_in_PopNB_mioi_oswt;
  assign accum_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff = accum_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp (
  clk, rst, act_in_PopNB_mioi_data_rsc_z_mxwt, act_in_PopNB_mioi_return_rsc_z_mxwt,
      act_in_PopNB_mioi_data_rsc_z, act_in_PopNB_mioi_biwt, act_in_PopNB_mioi_bdwt,
      act_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  output act_in_PopNB_mioi_return_rsc_z_mxwt;
  input [7:0] act_in_PopNB_mioi_data_rsc_z;
  input act_in_PopNB_mioi_biwt;
  input act_in_PopNB_mioi_bdwt;
  input act_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg act_in_PopNB_mioi_bcwt;
  reg [7:0] act_in_PopNB_mioi_data_rsc_z_bfwt;
  reg act_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign act_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_8_2_2(act_in_PopNB_mioi_data_rsc_z,
      act_in_PopNB_mioi_data_rsc_z_bfwt, act_in_PopNB_mioi_bcwt);
  assign act_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(act_in_PopNB_mioi_return_rsc_z,
      act_in_PopNB_mioi_return_rsc_z_bfwt, act_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_PopNB_mioi_bcwt <= 1'b0;
      act_in_PopNB_mioi_data_rsc_z_bfwt <= 8'b00000000;
      act_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      act_in_PopNB_mioi_bcwt <= ~((~(act_in_PopNB_mioi_bcwt | act_in_PopNB_mioi_biwt))
          | act_in_PopNB_mioi_bdwt);
      act_in_PopNB_mioi_data_rsc_z_bfwt <= act_in_PopNB_mioi_data_rsc_z_mxwt;
      act_in_PopNB_mioi_return_rsc_z_bfwt <= act_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl (
  PERun_wen, PERun_wten, act_in_PopNB_mioi_oswt, act_in_PopNB_mioi_biwt, act_in_PopNB_mioi_bdwt,
      act_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff, act_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input PERun_wten;
  input act_in_PopNB_mioi_oswt;
  output act_in_PopNB_mioi_biwt;
  output act_in_PopNB_mioi_bdwt;
  output act_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff;
  input act_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_PopNB_mioi_bdwt = act_in_PopNB_mioi_oswt & PERun_wen;
  assign act_in_PopNB_mioi_biwt = (~ PERun_wten) & act_in_PopNB_mioi_oswt;
  assign act_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff = act_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_out_PushNB_mioi_weight_out_PushNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_weight_out_PushNB_mioi_weight_out_PushNB_mio_wait_ctrl (
  PERun_wten, weight_out_PushNB_mioi_iswt0, weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct
);
  input PERun_wten;
  input weight_out_PushNB_mioi_iswt0;
  output weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;



  // Interconnect Declarations for Component Instantiations 
  assign weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct = weight_out_PushNB_mioi_iswt0
      & (~ PERun_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp (
  clk, rst, weight_in_PopNB_mioi_data_rsc_z_mxwt, weight_in_PopNB_mioi_return_rsc_z_mxwt,
      weight_in_PopNB_mioi_data_rsc_z, weight_in_PopNB_mioi_biwt, weight_in_PopNB_mioi_bdwt,
      weight_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  output weight_in_PopNB_mioi_return_rsc_z_mxwt;
  input [7:0] weight_in_PopNB_mioi_data_rsc_z;
  input weight_in_PopNB_mioi_biwt;
  input weight_in_PopNB_mioi_bdwt;
  input weight_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg weight_in_PopNB_mioi_bcwt;
  reg [7:0] weight_in_PopNB_mioi_data_rsc_z_bfwt;
  reg weight_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign weight_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_8_2_2(weight_in_PopNB_mioi_data_rsc_z,
      weight_in_PopNB_mioi_data_rsc_z_bfwt, weight_in_PopNB_mioi_bcwt);
  assign weight_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(weight_in_PopNB_mioi_return_rsc_z,
      weight_in_PopNB_mioi_return_rsc_z_bfwt, weight_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_in_PopNB_mioi_bcwt <= 1'b0;
      weight_in_PopNB_mioi_data_rsc_z_bfwt <= 8'b00000000;
      weight_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      weight_in_PopNB_mioi_bcwt <= ~((~(weight_in_PopNB_mioi_bcwt | weight_in_PopNB_mioi_biwt))
          | weight_in_PopNB_mioi_bdwt);
      weight_in_PopNB_mioi_data_rsc_z_bfwt <= weight_in_PopNB_mioi_data_rsc_z_mxwt;
      weight_in_PopNB_mioi_return_rsc_z_bfwt <= weight_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl (
  PERun_wen, weight_in_PopNB_mioi_oswt, PERun_wten, weight_in_PopNB_mioi_biwt, weight_in_PopNB_mioi_bdwt,
      weight_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff, weight_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input weight_in_PopNB_mioi_oswt;
  input PERun_wten;
  output weight_in_PopNB_mioi_biwt;
  output weight_in_PopNB_mioi_bdwt;
  output weight_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff;
  input weight_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign weight_in_PopNB_mioi_bdwt = weight_in_PopNB_mioi_oswt & PERun_wen;
  assign weight_in_PopNB_mioi_biwt = (~ PERun_wten) & weight_in_PopNB_mioi_oswt;
  assign weight_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff = weight_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi (
  clk, rst, accum_out_val, accum_out_rdy, accum_out_msg, PERun_wen, accum_out_Push_mioi_oswt,
      accum_out_Push_mioi_wen_comp, accum_out_Push_mioi_m_rsc_dat_PERun, accum_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;
  input PERun_wen;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_wen_comp;
  input [31:0] accum_out_Push_mioi_m_rsc_dat_PERun;
  input accum_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire accum_out_Push_mioi_biwt;
  wire accum_out_Push_mioi_bdwt;
  wire accum_out_Push_mioi_bcwt;
  wire accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  wire accum_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push  accum_out_Push_mioi
      (
      .this_val(accum_out_val),
      .this_rdy(accum_out_rdy),
      .this_msg(accum_out_msg),
      .m_rsc_dat(accum_out_Push_mioi_m_rsc_dat_PERun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .ccs_ccore_done_sync_vld(accum_out_Push_mioi_ccs_ccore_done_sync_vld)
    );
  SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .accum_out_Push_mioi_oswt(accum_out_Push_mioi_oswt),
      .accum_out_Push_mioi_biwt(accum_out_Push_mioi_biwt),
      .accum_out_Push_mioi_bdwt(accum_out_Push_mioi_bdwt),
      .accum_out_Push_mioi_bcwt(accum_out_Push_mioi_bcwt),
      .accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct(accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .accum_out_Push_mioi_ccs_ccore_done_sync_vld(accum_out_Push_mioi_ccs_ccore_done_sync_vld),
      .accum_out_Push_mioi_oswt_pff(accum_out_Push_mioi_oswt_pff)
    );
  SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .accum_out_Push_mioi_oswt(accum_out_Push_mioi_oswt),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_biwt(accum_out_Push_mioi_biwt),
      .accum_out_Push_mioi_bdwt(accum_out_Push_mioi_bdwt),
      .accum_out_Push_mioi_bcwt(accum_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi (
  clk, rst, act_out_val, act_out_rdy, act_out_msg, PERun_wen, act_out_Push_mioi_oswt,
      act_out_Push_mioi_wen_comp, act_out_Push_mioi_m_rsc_dat_PERun, act_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  input PERun_wen;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_wen_comp;
  input [7:0] act_out_Push_mioi_m_rsc_dat_PERun;
  input act_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_out_Push_mioi_biwt;
  wire act_out_Push_mioi_bdwt;
  wire act_out_Push_mioi_bcwt;
  wire act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  wire act_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_out_Push_mioi
      (
      .this_val(act_out_val),
      .this_rdy(act_out_rdy),
      .this_msg(act_out_msg),
      .m_rsc_dat(act_out_Push_mioi_m_rsc_dat_PERun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .ccs_ccore_done_sync_vld(act_out_Push_mioi_ccs_ccore_done_sync_vld)
    );
  SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .act_out_Push_mioi_oswt(act_out_Push_mioi_oswt),
      .act_out_Push_mioi_biwt(act_out_Push_mioi_biwt),
      .act_out_Push_mioi_bdwt(act_out_Push_mioi_bdwt),
      .act_out_Push_mioi_bcwt(act_out_Push_mioi_bcwt),
      .act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct(act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .act_out_Push_mioi_ccs_ccore_done_sync_vld(act_out_Push_mioi_ccs_ccore_done_sync_vld),
      .act_out_Push_mioi_oswt_pff(act_out_Push_mioi_oswt_pff)
    );
  SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_out_Push_mioi_oswt(act_out_Push_mioi_oswt),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .act_out_Push_mioi_biwt(act_out_Push_mioi_biwt),
      .act_out_Push_mioi_bdwt(act_out_Push_mioi_bdwt),
      .act_out_Push_mioi_bcwt(act_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi (
  clk, rst, accum_in_val, accum_in_rdy, accum_in_msg, PERun_wen, PERun_wten, accum_in_PopNB_mioi_oswt,
      accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_in_PopNB_mioi_return_rsc_z_mxwt,
      accum_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  input PERun_wen;
  input PERun_wten;
  input accum_in_PopNB_mioi_oswt;
  output [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  output accum_in_PopNB_mioi_return_rsc_z_mxwt;
  input accum_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [31:0] accum_in_PopNB_mioi_data_rsc_z;
  wire accum_in_PopNB_mioi_biwt;
  wire accum_in_PopNB_mioi_bdwt;
  wire accum_in_PopNB_mioi_return_rsc_z;
  wire accum_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB  accum_in_PopNB_mioi
      (
      .this_val(accum_in_val),
      .this_rdy(accum_in_rdy),
      .this_msg(accum_in_msg),
      .data_rsc_z(accum_in_PopNB_mioi_data_rsc_z),
      .do_wait_rsc_dat(accum_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff),
      .return_rsc_z(accum_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff)
    );
  SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .accum_in_PopNB_mioi_oswt(accum_in_PopNB_mioi_oswt),
      .accum_in_PopNB_mioi_biwt(accum_in_PopNB_mioi_biwt),
      .accum_in_PopNB_mioi_bdwt(accum_in_PopNB_mioi_bdwt),
      .accum_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff(accum_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff),
      .accum_in_PopNB_mioi_oswt_pff(accum_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .accum_in_PopNB_mioi_data_rsc_z_mxwt(accum_in_PopNB_mioi_data_rsc_z_mxwt),
      .accum_in_PopNB_mioi_return_rsc_z_mxwt(accum_in_PopNB_mioi_return_rsc_z_mxwt),
      .accum_in_PopNB_mioi_data_rsc_z(accum_in_PopNB_mioi_data_rsc_z),
      .accum_in_PopNB_mioi_biwt(accum_in_PopNB_mioi_biwt),
      .accum_in_PopNB_mioi_bdwt(accum_in_PopNB_mioi_bdwt),
      .accum_in_PopNB_mioi_return_rsc_z(accum_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi (
  clk, rst, act_in_val, act_in_rdy, act_in_msg, PERun_wen, PERun_wten, act_in_PopNB_mioi_oswt,
      act_in_PopNB_mioi_data_rsc_z_mxwt, act_in_PopNB_mioi_return_rsc_z_mxwt, act_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input PERun_wen;
  input PERun_wten;
  input act_in_PopNB_mioi_oswt;
  output [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  output act_in_PopNB_mioi_return_rsc_z_mxwt;
  input act_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [7:0] act_in_PopNB_mioi_data_rsc_z;
  wire act_in_PopNB_mioi_biwt;
  wire act_in_PopNB_mioi_bdwt;
  wire act_in_PopNB_mioi_return_rsc_z;
  wire act_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB  act_in_PopNB_mioi
      (
      .this_val(act_in_val),
      .this_rdy(act_in_rdy),
      .this_msg(act_in_msg),
      .data_rsc_z(act_in_PopNB_mioi_data_rsc_z),
      .do_wait_rsc_dat(act_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff),
      .return_rsc_z(act_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff)
    );
  SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_in_PopNB_mioi_oswt(act_in_PopNB_mioi_oswt),
      .act_in_PopNB_mioi_biwt(act_in_PopNB_mioi_biwt),
      .act_in_PopNB_mioi_bdwt(act_in_PopNB_mioi_bdwt),
      .act_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff(act_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff),
      .act_in_PopNB_mioi_oswt_pff(act_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_PopNB_mioi_data_rsc_z_mxwt(act_in_PopNB_mioi_data_rsc_z_mxwt),
      .act_in_PopNB_mioi_return_rsc_z_mxwt(act_in_PopNB_mioi_return_rsc_z_mxwt),
      .act_in_PopNB_mioi_data_rsc_z(act_in_PopNB_mioi_data_rsc_z),
      .act_in_PopNB_mioi_biwt(act_in_PopNB_mioi_biwt),
      .act_in_PopNB_mioi_bdwt(act_in_PopNB_mioi_bdwt),
      .act_in_PopNB_mioi_return_rsc_z(act_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_out_PushNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_weight_out_PushNB_mioi (
  clk, rst, weight_out_val, weight_out_rdy, weight_out_msg, PERun_wten, weight_out_PushNB_mioi_iswt0,
      weight_out_PushNB_mioi_m_rsc_dat_PERun
);
  input clk;
  input rst;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;
  input PERun_wten;
  input weight_out_PushNB_mioi_iswt0;
  input [7:0] weight_out_PushNB_mioi_m_rsc_dat_PERun;


  // Interconnect Declarations
  wire weight_out_PushNB_mioi_return_rsc_z;
  wire weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB  weight_out_PushNB_mioi
      (
      .this_val(weight_out_val),
      .this_rdy(weight_out_rdy),
      .this_msg(weight_out_msg),
      .m_rsc_dat(weight_out_PushNB_mioi_m_rsc_dat_PERun),
      .return_rsc_z(weight_out_PushNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
  SysPE_PERun_weight_out_PushNB_mioi_weight_out_PushNB_mio_wait_ctrl SysPE_PERun_weight_out_PushNB_mioi_weight_out_PushNB_mio_wait_ctrl_inst
      (
      .PERun_wten(PERun_wten),
      .weight_out_PushNB_mioi_iswt0(weight_out_PushNB_mioi_iswt0),
      .weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct(weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, PERun_wen, weight_in_PopNB_mioi_oswt,
      PERun_wten, weight_in_PopNB_mioi_data_rsc_z_mxwt, weight_in_PopNB_mioi_return_rsc_z_mxwt,
      weight_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input PERun_wen;
  input weight_in_PopNB_mioi_oswt;
  input PERun_wten;
  output [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  output weight_in_PopNB_mioi_return_rsc_z_mxwt;
  input weight_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [7:0] weight_in_PopNB_mioi_data_rsc_z;
  wire weight_in_PopNB_mioi_biwt;
  wire weight_in_PopNB_mioi_bdwt;
  wire weight_in_PopNB_mioi_return_rsc_z;
  wire weight_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_in_PopNB_mioi
      (
      .this_val(weight_in_val),
      .this_rdy(weight_in_rdy),
      .this_msg(weight_in_msg),
      .data_rsc_z(weight_in_PopNB_mioi_data_rsc_z),
      .do_wait_rsc_dat(weight_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff),
      .return_rsc_z(weight_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff)
    );
  SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .weight_in_PopNB_mioi_oswt(weight_in_PopNB_mioi_oswt),
      .PERun_wten(PERun_wten),
      .weight_in_PopNB_mioi_biwt(weight_in_PopNB_mioi_biwt),
      .weight_in_PopNB_mioi_bdwt(weight_in_PopNB_mioi_bdwt),
      .weight_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_pff(weight_in_PopNB_mioi_do_wait_rsc_dat_PERun_sct_iff),
      .weight_in_PopNB_mioi_oswt_pff(weight_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .weight_in_PopNB_mioi_data_rsc_z_mxwt(weight_in_PopNB_mioi_data_rsc_z_mxwt),
      .weight_in_PopNB_mioi_return_rsc_z_mxwt(weight_in_PopNB_mioi_return_rsc_z_mxwt),
      .weight_in_PopNB_mioi_data_rsc_z(weight_in_PopNB_mioi_data_rsc_z),
      .weight_in_PopNB_mioi_biwt(weight_in_PopNB_mioi_biwt),
      .weight_in_PopNB_mioi_bdwt(weight_in_PopNB_mioi_bdwt),
      .weight_in_PopNB_mioi_return_rsc_z(weight_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun
// ------------------------------------------------------------------


module SysPE_PERun (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, act_in_val, act_in_rdy,
      act_in_msg, accum_in_val, accum_in_rdy, accum_in_msg, act_out_val, act_out_rdy,
      act_out_msg, accum_out_val, accum_out_rdy, accum_out_msg, weight_out_val, weight_out_rdy,
      weight_out_msg
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;


  // Interconnect Declarations
  wire PERun_wen;
  wire PERun_wten;
  wire [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  wire weight_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  wire act_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  wire accum_in_PopNB_mioi_return_rsc_z_mxwt;
  wire act_out_Push_mioi_wen_comp;
  wire accum_out_Push_mioi_wen_comp;
  wire [1:0] fsm_output;
  wire while_while_or_tmp;
  wire is_accum_in_sva_dfm_1;
  reg is_accum_in_sva;
  reg while_stage_0_3;
  reg is_act_in_sva;
  wire while_land_lpi_1_dfm_1;
  reg reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  wire is_accum_in_and_cse;
  wire and_1_cse;
  wire and_5_rmff;
  wire and_4_rmff;
  reg [7:0] act_reg_sva;
  wire [7:0] act_out_Push_mioi_m_rsc_dat_PERun_mx1;
  reg [7:0] weight_reg_sva;
  wire [31:0] accum_reg_sva_mx0;
  reg [31:0] accum_reg_sva;

  wire[0:0] mux_7_nl;
  wire[0:0] or_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_11_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] nor_1_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] nor_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff;
  assign nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff =
      fsm_output[1];
  wire [0:0] nl_SysPE_PERun_weight_out_PushNB_mioi_inst_PERun_wten;
  assign nl_SysPE_PERun_weight_out_PushNB_mioi_inst_PERun_wten = ~ PERun_wen;
  wire [0:0] nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_iswt0;
  assign nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_iswt0
      = reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse & weight_in_PopNB_mioi_return_rsc_z_mxwt;
  wire[0:0] or_nl;
  wire [7:0] nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun;
  assign or_nl = is_act_in_sva | (fsm_output[0]);
  assign nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun
      = MUX_v_8_2_2(act_in_PopNB_mioi_data_rsc_z_mxwt, act_reg_sva, or_nl);
  wire[15:0] while_if_3_accum_out_reg_mul_nl;
  wire [31:0] nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun;
  assign while_if_3_accum_out_reg_mul_nl = conv_s2u_16_16($signed((act_out_Push_mioi_m_rsc_dat_PERun_mx1))
      * $signed(weight_reg_sva));
  assign nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun
      = conv_s2u_16_32(while_if_3_accum_out_reg_mul_nl) + accum_reg_sva_mx0;
  SysPE_PERun_weight_in_PopNB_mioi SysPE_PERun_weight_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_val),
      .weight_in_rdy(weight_in_rdy),
      .weight_in_msg(weight_in_msg),
      .PERun_wen(PERun_wen),
      .weight_in_PopNB_mioi_oswt(reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .PERun_wten(PERun_wten),
      .weight_in_PopNB_mioi_data_rsc_z_mxwt(weight_in_PopNB_mioi_data_rsc_z_mxwt),
      .weight_in_PopNB_mioi_return_rsc_z_mxwt(weight_in_PopNB_mioi_return_rsc_z_mxwt),
      .weight_in_PopNB_mioi_oswt_pff(nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff[0:0])
    );
  SysPE_PERun_weight_out_PushNB_mioi SysPE_PERun_weight_out_PushNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .weight_out_val(weight_out_val),
      .weight_out_rdy(weight_out_rdy),
      .weight_out_msg(weight_out_msg),
      .PERun_wten(nl_SysPE_PERun_weight_out_PushNB_mioi_inst_PERun_wten[0:0]),
      .weight_out_PushNB_mioi_iswt0(nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_iswt0[0:0]),
      .weight_out_PushNB_mioi_m_rsc_dat_PERun(weight_in_PopNB_mioi_data_rsc_z_mxwt)
    );
  SysPE_PERun_act_in_PopNB_mioi SysPE_PERun_act_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .act_in_val(act_in_val),
      .act_in_rdy(act_in_rdy),
      .act_in_msg(act_in_msg),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_in_PopNB_mioi_oswt(reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .act_in_PopNB_mioi_data_rsc_z_mxwt(act_in_PopNB_mioi_data_rsc_z_mxwt),
      .act_in_PopNB_mioi_return_rsc_z_mxwt(act_in_PopNB_mioi_return_rsc_z_mxwt),
      .act_in_PopNB_mioi_oswt_pff(and_5_rmff)
    );
  SysPE_PERun_accum_in_PopNB_mioi SysPE_PERun_accum_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .accum_in_val(accum_in_val),
      .accum_in_rdy(accum_in_rdy),
      .accum_in_msg(accum_in_msg),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .accum_in_PopNB_mioi_oswt(reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .accum_in_PopNB_mioi_data_rsc_z_mxwt(accum_in_PopNB_mioi_data_rsc_z_mxwt),
      .accum_in_PopNB_mioi_return_rsc_z_mxwt(accum_in_PopNB_mioi_return_rsc_z_mxwt),
      .accum_in_PopNB_mioi_oswt_pff(and_4_rmff)
    );
  SysPE_PERun_act_out_Push_mioi SysPE_PERun_act_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .act_out_val(act_out_val),
      .act_out_rdy(act_out_rdy),
      .act_out_msg(act_out_msg),
      .PERun_wen(PERun_wen),
      .act_out_Push_mioi_oswt(reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .act_out_Push_mioi_m_rsc_dat_PERun(nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun[7:0]),
      .act_out_Push_mioi_oswt_pff(and_1_cse)
    );
  SysPE_PERun_accum_out_Push_mioi SysPE_PERun_accum_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .accum_out_val(accum_out_val),
      .accum_out_rdy(accum_out_rdy),
      .accum_out_msg(accum_out_msg),
      .PERun_wen(PERun_wen),
      .accum_out_Push_mioi_oswt(reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_m_rsc_dat_PERun(nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun[31:0]),
      .accum_out_Push_mioi_oswt_pff(and_1_cse)
    );
  SysPE_PERun_staller SysPE_PERun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp)
    );
  SysPE_PERun_PERun_fsm SysPE_PERun_PERun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PERun_wen(PERun_wen),
      .fsm_output(fsm_output)
    );
  assign and_1_cse = while_while_or_tmp & is_accum_in_sva_dfm_1 & while_stage_0_3;
  assign or_9_nl = (~ is_accum_in_sva_dfm_1) | act_in_PopNB_mioi_return_rsc_z_mxwt
      | is_act_in_sva;
  assign mux_7_nl = MUX_s_1_2_2((~ is_accum_in_sva), (or_9_nl), while_stage_0_3);
  assign and_4_rmff = (mux_7_nl) & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  assign or_11_nl = is_accum_in_sva_dfm_1 | (~ while_while_or_tmp);
  assign mux_8_nl = MUX_s_1_2_2((~ is_act_in_sva), (or_11_nl), while_stage_0_3);
  assign and_5_rmff = (mux_8_nl) & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  assign is_accum_in_and_cse = PERun_wen & while_stage_0_3;
  assign act_out_Push_mioi_m_rsc_dat_PERun_mx1 = MUX_v_8_2_2(act_in_PopNB_mioi_data_rsc_z_mxwt,
      act_reg_sva, is_act_in_sva);
  assign accum_reg_sva_mx0 = MUX_v_32_2_2(accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_reg_sva,
      is_accum_in_sva);
  assign is_accum_in_sva_dfm_1 = accum_in_PopNB_mioi_return_rsc_z_mxwt | is_accum_in_sva;
  assign while_land_lpi_1_dfm_1 = is_accum_in_sva_dfm_1 & while_while_or_tmp;
  assign while_while_or_tmp = act_in_PopNB_mioi_return_rsc_z_mxwt | is_act_in_sva;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      while_stage_0_3 <= 1'b0;
    end
    else if ( PERun_wen ) begin
      reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_1_cse;
      reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_4_rmff;
      reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_5_rmff;
      reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= fsm_output[1];
      while_stage_0_3 <= reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      is_accum_in_sva <= 1'b0;
      is_act_in_sva <= 1'b0;
    end
    else if ( is_accum_in_and_cse ) begin
      is_accum_in_sva <= is_accum_in_sva_dfm_1 & (~ while_land_lpi_1_dfm_1);
      is_act_in_sva <= while_while_or_tmp & (~ while_land_lpi_1_dfm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_reg_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( PERun_wen & (mux_5_nl) ) begin
      accum_reg_sva <= accum_reg_sva_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_reg_sva <= 8'b00000000;
    end
    else if ( PERun_wen & (mux_6_nl) ) begin
      act_reg_sva <= act_out_Push_mioi_m_rsc_dat_PERun_mx1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_reg_sva <= 8'b00000000;
    end
    else if ( PERun_wen & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse
        & weight_in_PopNB_mioi_return_rsc_z_mxwt ) begin
      weight_reg_sva <= weight_in_PopNB_mioi_data_rsc_z_mxwt;
    end
  end
  assign nor_1_nl = ~((~ is_accum_in_sva_dfm_1) | act_in_PopNB_mioi_return_rsc_z_mxwt
      | is_act_in_sva);
  assign mux_5_nl = MUX_s_1_2_2(is_accum_in_sva, (nor_1_nl), while_stage_0_3);
  assign nor_nl = ~(is_accum_in_sva_dfm_1 | (~ while_while_or_tmp));
  assign mux_6_nl = MUX_s_1_2_2(is_act_in_sva, (nor_nl), while_stage_0_3);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [15:0] conv_s2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_16 = vector;
  end
  endfunction


  function automatic [31:0] conv_s2u_16_32 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_32 = {{16{vector[15]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_rtl
// ------------------------------------------------------------------


module SysPE_rtl (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, act_in_val, act_in_rdy,
      act_in_msg, accum_in_val, accum_in_rdy, accum_in_msg, act_out_val, act_out_rdy,
      act_out_msg, accum_out_val, accum_out_rdy, accum_out_msg, weight_out_val, weight_out_rdy,
      weight_out_msg
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;



  // Interconnect Declarations for Component Instantiations 
  SysPE_PERun SysPE_PERun_inst (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_val),
      .weight_in_rdy(weight_in_rdy),
      .weight_in_msg(weight_in_msg),
      .act_in_val(act_in_val),
      .act_in_rdy(act_in_rdy),
      .act_in_msg(act_in_msg),
      .accum_in_val(accum_in_val),
      .accum_in_rdy(accum_in_rdy),
      .accum_in_msg(accum_in_msg),
      .act_out_val(act_out_val),
      .act_out_rdy(act_out_rdy),
      .act_out_msg(act_out_msg),
      .accum_out_val(accum_out_val),
      .accum_out_rdy(accum_out_rdy),
      .accum_out_msg(accum_out_msg),
      .weight_out_val(weight_out_val),
      .weight_out_rdy(weight_out_rdy),
      .weight_out_msg(weight_out_msg)
    );
endmodule



