
//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_out_dreg_v2.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module mgc_out_dreg_v2 (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_in_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2017 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------


module ccs_in_v1 (idat, dat);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] idat;
  input  [width-1:0] dat;

  wire   [width-1:0] idat;

  assign idat = dat;

endmodule


//------> ../td_ccore_solutions/Connections__Combinational_ArbitratedScratchpad_InputSetup--_31ec8cab963b6f5e97b0c13f1550d1c18e15_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:10:20 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PopNB_core
    (
  this_val, this_rdy, this_msg, data_type_val_rsc_z, data_valids_rsc_z, data_addr_rsc_z,
      data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [136:0] this_msg;
  output data_type_val_rsc_z;
  output [7:0] data_valids_rsc_z;
  output [63:0] data_addr_rsc_z;
  output [63:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_data_type_val_rsci_d;
  assign nl_data_type_val_rsci_d = this_msg[136];
  wire [7:0] nl_data_valids_rsci_d;
  assign nl_data_valids_rsci_d = {(this_msg[135]) , (this_msg[118]) , (this_msg[101])
      , (this_msg[84]) , (this_msg[67]) , (this_msg[50]) , (this_msg[33]) , (this_msg[16])};
  wire [63:0] nl_data_addr_rsci_d;
  assign nl_data_addr_rsci_d = {(this_msg[134:127]) , (this_msg[117:110]) , (this_msg[100:93])
      , (this_msg[83:76]) , (this_msg[66:59]) , (this_msg[49:42]) , (this_msg[32:25])
      , (this_msg[15:8])};
  wire [63:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = {(this_msg[126:119]) , (this_msg[109:102]) , (this_msg[92:85])
      , (this_msg[75:68]) , (this_msg[58:51]) , (this_msg[41:34]) , (this_msg[24:17])
      , (this_msg[7:0])};
  mgc_out_dreg_v2 #(.rscid(32'sd215),
  .width(32'sd1)) data_type_val_rsci (
      .d(nl_data_type_val_rsci_d[0:0]),
      .z(data_type_val_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd216),
  .width(32'sd8)) data_valids_rsci (
      .d(nl_data_valids_rsci_d[7:0]),
      .z(data_valids_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd217),
  .width(32'sd64)) data_addr_rsci (
      .d(nl_data_addr_rsci_d[63:0]),
      .z(data_addr_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd218),
  .width(32'sd64)) data_data_rsci (
      .d(nl_data_data_rsci_d[63:0]),
      .z(data_data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd219),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd322),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PopNB
    (
  this_val, this_rdy, this_msg, data_type_val_rsc_z, data_valids_rsc_z, data_addr_rsc_z,
      data_data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [136:0] this_msg;
  output data_type_val_rsc_z;
  output [7:0] data_valids_rsc_z;
  output [63:0] data_addr_rsc_z;
  output [63:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PopNB_core
      Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_type_val_rsc_z(data_type_val_rsc_z),
      .data_valids_rsc_z(data_valids_rsc_z),
      .data_addr_rsc_z(data_addr_rsc_z),
      .data_data_rsc_z(data_data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__InBlocking_InputSetup__WriteReq_Connections__--_749f9cf99c5bf2b4f3e6a99e1ab903e16fa4_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:10:16 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_InputSetup_WriteReq_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_InBlocking_InputSetup_WriteReq_Connections_SYN_PORT_PopNB_core
    (
  this_val, this_rdy, this_msg, data_data_data_rsc_z, data_index_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [68:0] this_msg;
  output [63:0] data_data_data_rsc_z;
  output [4:0] data_index_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_data_data_data_rsci_d;
  assign nl_data_data_data_rsci_d = this_msg[63:0];
  wire [4:0] nl_data_index_rsci_d;
  assign nl_data_index_rsci_d = this_msg[68:64];
  mgc_out_dreg_v2 #(.rscid(32'sd223),
  .width(32'sd64)) data_data_data_rsci (
      .d(nl_data_data_data_rsci_d[63:0]),
      .z(data_data_data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd224),
  .width(32'sd5)) data_index_rsci (
      .d(nl_data_index_rsci_d[4:0]),
      .z(data_index_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd226),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd321),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_InputSetup_WriteReq_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_InBlocking_InputSetup_WriteReq_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_data_data_rsc_z, data_index_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [68:0] this_msg;
  output [63:0] data_data_data_rsc_z;
  output [4:0] data_index_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_InputSetup_WriteReq_Connections_SYN_PORT_PopNB_core Connections_InBlocking_InputSetup_WriteReq_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_data_data_rsc_z(data_data_data_rsc_z),
      .data_index_rsc_z(data_index_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ccs_sync_out_vld_v1.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ccs_sync_out_vld_v1 (vld, ivld);
  parameter integer rscid = 1;

  input  ivld;
  output vld;

  wire   vld;

  assign vld = ivld;
endmodule

//------> ../td_ccore_solutions/Connections__Combinational_ArbitratedScratchpad_InputSetup--_6d01a7417bfbe5463c65573f0d893d1a73e5_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:10:12 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_Push_core
    (
  this_val, this_rdy, this_msg, m_valids_rsc_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [71:0] this_msg;
  input [7:0] m_valids_rsc_dat;
  input [63:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [7:0] m_valids_rsci_idat;
  wire [63:0] m_data_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg wm_val_Marshall_72U_for_8_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_72U_for_8_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1;
  reg wm_val_Marshall_72U_for_7_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_72U_for_7_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1;
  reg wm_val_Marshall_72U_for_6_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_72U_for_6_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1;
  reg wm_val_Marshall_72U_for_5_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_72U_for_5_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1;
  reg wm_val_Marshall_72U_for_4_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_72U_for_4_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1;
  reg wm_val_Marshall_72U_for_3_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_72U_for_3_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1;
  reg wm_val_Marshall_72U_for_2_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_72U_for_2_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1;
  reg wm_val_Marshall_72U_for_1_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_72U_for_1_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_2;
  wire and_dcpl_5;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire and_cse;
  wire or_5_cse;
  reg [7:0] m_valids_buf_lpi_1_dfm;
  reg [63:0] m_data_buf_lpi_1_dfm;
  wire this_val_mx0c1;
  wire [7:0] m_valids_buf_lpi_1_dfm_mx0;
  wire [63:0] m_data_buf_lpi_1_dfm_mx0;
  wire and_6_cse;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd228),
  .width(32'sd8)) m_valids_rsci (
      .dat(m_valids_rsc_dat),
      .idat(m_valids_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd229),
  .width(32'sd64)) m_data_rsci (
      .dat(m_data_rsc_dat),
      .idat(m_data_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd320),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd331)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign this_msg = {wm_val_Marshall_72U_for_8_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_72U_for_8_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
      , wm_val_Marshall_72U_for_7_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_72U_for_7_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
      , wm_val_Marshall_72U_for_6_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_72U_for_6_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
      , wm_val_Marshall_72U_for_5_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_72U_for_5_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
      , wm_val_Marshall_72U_for_4_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_72U_for_4_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
      , wm_val_Marshall_72U_for_3_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_72U_for_3_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
      , wm_val_Marshall_72U_for_2_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_72U_for_2_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
      , wm_val_Marshall_72U_for_1_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_72U_for_1_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_2};
  assign and_6_cse = (this_rdy | (~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1))
      & ccs_ccore_start_rsci_idat;
  assign or_5_cse = ccs_ccore_start_rsci_idat | and_cse;
  assign m_valids_buf_lpi_1_dfm_mx0 = MUX_v_8_2_2(m_valids_rsci_idat, m_valids_buf_lpi_1_dfm,
      and_cse);
  assign m_data_buf_lpi_1_dfm_mx0 = MUX_v_64_2_2(m_data_rsci_idat, m_data_buf_lpi_1_dfm,
      and_cse);
  assign and_cse = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign and_dcpl_5 = ~((~((~ io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1) | this_rdy))
      | ccs_ccore_start_rsci_idat);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_5_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_8_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_8_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_buf_lpi_1_dfm_mx0[7];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_8_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= 8'b00000000;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_8_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= m_data_buf_lpi_1_dfm_mx0[63:56];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_7_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_7_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_buf_lpi_1_dfm_mx0[6];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_7_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= 8'b00000000;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_7_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= m_data_buf_lpi_1_dfm_mx0[55:48];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_6_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_6_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_buf_lpi_1_dfm_mx0[5];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_6_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= 8'b00000000;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_6_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= m_data_buf_lpi_1_dfm_mx0[47:40];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_5_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_5_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_buf_lpi_1_dfm_mx0[4];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_5_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= 8'b00000000;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_5_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= m_data_buf_lpi_1_dfm_mx0[39:32];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_4_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_4_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_buf_lpi_1_dfm_mx0[3];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_4_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= 8'b00000000;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_4_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= m_data_buf_lpi_1_dfm_mx0[31:24];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_3_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_3_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_buf_lpi_1_dfm_mx0[2];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_3_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= 8'b00000000;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_3_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= m_data_buf_lpi_1_dfm_mx0[23:16];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_2_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_2_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_buf_lpi_1_dfm_mx0[1];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_2_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= 8'b00000000;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_2_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_1
          <= m_data_buf_lpi_1_dfm_mx0[15:8];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_1_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_1_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_buf_lpi_1_dfm_mx0[0];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_72U_for_1_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_2
          <= 8'b00000000;
    end
    else if ( ~ and_dcpl_5 ) begin
      wm_val_Marshall_72U_for_1_to_sc_8_v_slc_this_write_msg_wm_val_data_8_7_0_2
          <= m_data_buf_lpi_1_dfm_mx0[7:0];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      m_valids_buf_lpi_1_dfm <= 8'b00000000;
      m_data_buf_lpi_1_dfm <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( and_6_cse ) begin
      m_valids_buf_lpi_1_dfm <= m_valids_buf_lpi_1_dfm_mx0;
      m_data_buf_lpi_1_dfm <= m_data_buf_lpi_1_dfm_mx0;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_5_cse;
    end
  end

  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_Push
    (
  this_val, this_rdy, this_msg, m_valids_rsc_dat, m_data_rsc_dat, ccs_ccore_start_rsc_dat,
      ccs_ccore_done_sync_vld, ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [71:0] this_msg;
  input [7:0] m_valids_rsc_dat;
  input [63:0] m_data_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_Push_core
      Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_valids_rsc_dat(m_valids_rsc_dat),
      .m_data_rsc_dat(m_data_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/mgc_shift_l_beh_v5.v 
module mgc_shift_l_v5(a,s,z);
   parameter    width_a = 4;
   parameter    signd_a = 1;
   parameter    width_s = 2;
   parameter    width_z = 8;

   input [width_a-1:0] a;
   input [width_s-1:0] s;
   output [width_z -1:0] z;

   generate
   if (signd_a)
   begin: SGNED
      assign z = fshl_u(a,s,a[width_a-1]);
   end
   else
   begin: UNSGNED
      assign z = fshl_u(a,s,1'b0);
   end
   endgenerate

   //Shift-left - unsigned shift argument one bit more
   function [width_z-1:0] fshl_u_1;
      input [width_a  :0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      parameter olen = width_z;
      parameter ilen = width_a+1;
      parameter len = (ilen >= olen) ? ilen : olen;
      reg [len-1:0] result;
      reg [len-1:0] result_t;
      begin
        result_t = {(len){sbit}};
        result_t[ilen-1:0] = arg1;
        result = result_t <<< arg2;
        fshl_u_1 =  result[olen-1:0];
      end
   endfunction // fshl_u

   //Shift-left - unsigned shift argument
   function [width_z-1:0] fshl_u;
      input [width_a-1:0] arg1;
      input [width_s-1:0] arg2;
      input sbit;
      fshl_u = fshl_u_1({sbit,arg1} ,arg2, sbit);
   endfunction // fshl_u

endmodule

//------> ../td_ccore_solutions/Connections__InBlocking_InputSetup__StartType_Connections_--_5b702d3f41a65f0c5ddd48c1b46b684e599a_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:10:07 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_InputSetup_StartType_Connections_SYN_PORT_Pop_core
// ------------------------------------------------------------------


module Connections_InBlocking_InputSetup_StartType_Connections_SYN_PORT_Pop_core
    (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [5:0] this_msg;
  output [5:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_2_cse;
  wire this_rdy_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [5:0] nl_return_rsci_d;
  assign nl_return_rsci_d = this_msg;
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_val;
  mgc_out_dreg_v2 #(.rscid(32'sd232),
  .width(32'sd6)) return_rsci (
      .d(nl_return_rsci_d[5:0]),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd319),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd330)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_2_cse = ccs_ccore_start_rsci_idat | (io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & (~ this_val));
  assign this_rdy_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_val
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( or_2_cse | this_rdy_mx0c1 ) begin
      this_rdy <= ~ this_rdy_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_2_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_InputSetup_StartType_Connections_SYN_PORT_Pop
// ------------------------------------------------------------------


module Connections_InBlocking_InputSetup_StartType_Connections_SYN_PORT_Pop (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [5:0] this_msg;
  output [5:0] return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_InputSetup_StartType_Connections_SYN_PORT_Pop_core Connections_InBlocking_InputSetup_StartType_Connections_SYN_PORT_Pop_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_ArbitratedScratchpad_InputSetup--_694dcb83f2aefc5cd19d731ef7b159598485_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:10:03 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PushNB_core
// ------------------------------------------------------------------


module Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PushNB_core
    (
  this_val, this_rdy, this_msg, m_valids_rsc_dat, m_addr_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [136:0] this_msg;
  input [7:0] m_valids_rsc_dat;
  input [63:0] m_addr_rsc_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [7:0] m_valids_rsci_idat;
  wire [63:0] m_addr_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  reg wm_val_Marshall_137U_for_8_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_137U_for_8_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1;
  reg wm_val_Marshall_137U_for_7_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_137U_for_7_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1;
  reg wm_val_Marshall_137U_for_6_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_137U_for_6_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1;
  reg wm_val_Marshall_137U_for_5_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_137U_for_5_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1;
  reg wm_val_Marshall_137U_for_4_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_137U_for_4_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1;
  reg wm_val_Marshall_137U_for_3_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_137U_for_3_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1;
  reg wm_val_Marshall_137U_for_2_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_137U_for_2_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1;
  reg wm_val_Marshall_137U_for_1_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1;
  reg [7:0] wm_val_Marshall_137U_for_1_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd234),
  .width(32'sd8)) m_valids_rsci (
      .dat(m_valids_rsc_dat),
      .idat(m_valids_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd235),
  .width(32'sd64)) m_addr_rsci (
      .dat(m_addr_rsc_dat),
      .idat(m_addr_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd237),
  .width(32'sd1)) return_rsci (
      .d(this_rdy),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd318),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign this_msg = {1'b0 , wm_val_Marshall_137U_for_8_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_137U_for_8_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
      , 8'b00000000 , wm_val_Marshall_137U_for_7_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_137U_for_7_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
      , 8'b00000000 , wm_val_Marshall_137U_for_6_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_137U_for_6_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
      , 8'b00000000 , wm_val_Marshall_137U_for_5_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_137U_for_5_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
      , 8'b00000000 , wm_val_Marshall_137U_for_4_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_137U_for_4_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
      , 8'b00000000 , wm_val_Marshall_137U_for_3_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_137U_for_3_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
      , 8'b00000000 , wm_val_Marshall_137U_for_2_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_137U_for_2_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
      , 8'b00000000 , wm_val_Marshall_137U_for_1_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
      , wm_val_Marshall_137U_for_1_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
      , 8'b00000000};
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_val <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      wm_val_Marshall_137U_for_8_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
      wm_val_Marshall_137U_for_8_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= 8'b00000000;
      wm_val_Marshall_137U_for_7_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
      wm_val_Marshall_137U_for_7_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= 8'b00000000;
      wm_val_Marshall_137U_for_6_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
      wm_val_Marshall_137U_for_6_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= 8'b00000000;
      wm_val_Marshall_137U_for_5_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
      wm_val_Marshall_137U_for_5_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= 8'b00000000;
      wm_val_Marshall_137U_for_4_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
      wm_val_Marshall_137U_for_4_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= 8'b00000000;
      wm_val_Marshall_137U_for_3_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
      wm_val_Marshall_137U_for_3_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= 8'b00000000;
      wm_val_Marshall_137U_for_2_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
      wm_val_Marshall_137U_for_2_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= 8'b00000000;
      wm_val_Marshall_137U_for_1_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= 1'b0;
      wm_val_Marshall_137U_for_1_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= 8'b00000000;
    end
    else if ( ccs_ccore_start_rsci_idat ) begin
      wm_val_Marshall_137U_for_8_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_rsci_idat[7];
      wm_val_Marshall_137U_for_8_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= m_addr_rsci_idat[63:56];
      wm_val_Marshall_137U_for_7_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_rsci_idat[6];
      wm_val_Marshall_137U_for_7_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= m_addr_rsci_idat[55:48];
      wm_val_Marshall_137U_for_6_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_rsci_idat[5];
      wm_val_Marshall_137U_for_6_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= m_addr_rsci_idat[47:40];
      wm_val_Marshall_137U_for_5_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_rsci_idat[4];
      wm_val_Marshall_137U_for_5_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= m_addr_rsci_idat[39:32];
      wm_val_Marshall_137U_for_4_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_rsci_idat[3];
      wm_val_Marshall_137U_for_4_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= m_addr_rsci_idat[31:24];
      wm_val_Marshall_137U_for_3_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_rsci_idat[2];
      wm_val_Marshall_137U_for_3_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= m_addr_rsci_idat[23:16];
      wm_val_Marshall_137U_for_2_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_rsci_idat[1];
      wm_val_Marshall_137U_for_2_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= m_addr_rsci_idat[15:8];
      wm_val_Marshall_137U_for_1_type_to_vector_bool_1_slc_this_write_msg_wm_val_valids_1_0_1
          <= m_valids_rsci_idat[0];
      wm_val_Marshall_137U_for_1_to_sc_8_1_v_slc_this_write_msg_wm_val_addr_8_7_0_1
          <= m_addr_rsci_idat[7:0];
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PushNB
// ------------------------------------------------------------------


module Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PushNB
    (
  this_val, this_rdy, this_msg, m_valids_rsc_dat, m_addr_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [136:0] this_msg;
  input [7:0] m_valids_rsc_dat;
  input [63:0] m_addr_rsc_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PushNB_core
      Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PushNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_valids_rsc_dat(m_valids_rsc_dat),
      .m_addr_rsc_dat(m_addr_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_ArbitratedScratchpad_InputSetup--_a25023c05ca59912d81479e03633279876b3_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:09:59 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_PopNB_core
    (
  this_val, this_rdy, this_msg, data_valids_rsc_z, data_data_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [71:0] this_msg;
  output [7:0] data_valids_rsc_z;
  output [63:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_data_valids_rsci_d;
  assign nl_data_valids_rsci_d = {(this_msg[71]) , (this_msg[62]) , (this_msg[53])
      , (this_msg[44]) , (this_msg[35]) , (this_msg[26]) , (this_msg[17]) , (this_msg[8])};
  wire [63:0] nl_data_data_rsci_d;
  assign nl_data_data_rsci_d = {(this_msg[70:63]) , (this_msg[61:54]) , (this_msg[52:45])
      , (this_msg[43:36]) , (this_msg[34:27]) , (this_msg[25:18]) , (this_msg[16:9])
      , (this_msg[7:0])};
  mgc_out_dreg_v2 #(.rscid(32'sd241),
  .width(32'sd8)) data_valids_rsci (
      .d(nl_data_valids_rsci_d[7:0]),
      .z(data_valids_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd242),
  .width(32'sd64)) data_data_rsci (
      .d(nl_data_data_rsci_d[63:0]),
      .z(data_data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd243),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd317),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_PopNB
    (
  this_val, this_rdy, this_msg, data_valids_rsc_z, data_data_rsc_z, return_rsc_z,
      ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [71:0] this_msg;
  output [7:0] data_valids_rsc_z;
  output [63:0] data_data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_PopNB_core
      Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_valids_rsc_z(data_valids_rsc_z),
      .data_data_rsc_z(data_data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__OutBlocking_SysPE__InputType_Connections__SYN--_0915a3f7c0fd3ff66acab9cdc0d4268d5eed_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:09:42 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [7:0] this_msg;
  reg [7:0] this_msg;
  input [7:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [7:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd10),
  .width(32'sd8)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd326),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd333)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 8'b00000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_msg <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [7:0] this_msg;
  input [7:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> /cad/tools/mentor/catapult/Catapult_Synthesis_10.4b-841621/Mgc_home/pkgs/siflibs/ram_sync_single_be_generic.v 
//------------------------------------------------------------------------------
// Catapult Synthesis - Sample I/O Port Library
//
// Copyright (c) 2003-2015 Mentor Graphics Corp.
//       All Rights Reserved
//
// This document may be used and distributed without restriction provided that
// this copyright statement is not removed from the file and that any derivative
// work contains this copyright notice.
//
// The design information contained in this file is intended to be an example
// of the functionality which the end user may study in preparation for creating
// their own custom interfaces. This design does not necessarily present a 
// complete implementation of the named protocol or standard.
//
//------------------------------------------------------------------------------

module ram_sync_single_be ( data_in, addr, re, we, data_out, clk, a_rst, s_rst, en);

  parameter ram_id = 1;
  parameter words = 'd16;
  parameter width = 'd16;
  parameter addr_width = 4;
  parameter [0:0] a_reset_active = 1;
  parameter [0:0] s_reset_active = 1;
  parameter [0:0] enable_active = 1;
  parameter [0:0] re_active = 1;
  parameter [0:0] we_active = 1;
  parameter num_byte_enables = 1;
  parameter [0:0] clock_edge = 1;
  parameter no_of_RAM_readwrite_port = 1;

  localparam byte_width = width / num_byte_enables;


  input [width-1:0] data_in;
  input [addr_width-1:0] addr;
  input [num_byte_enables-1:0] re;
  input [num_byte_enables-1:0] we;
  output reg [width-1:0] data_out;
  input clk;
  input a_rst;
  input s_rst;
  input en;

  // synopsys translate_off
  reg  [addr_width-1:0] addr_reg;
  reg  [num_byte_enables-1:0] re_reg;
  reg  [width-1:0] mem [words-1:0];  

  integer count;
  initial
  begin
    for (count = 0; count < words; count = count + 1)
      mem[count] = 0;
  end

  integer i;
  generate
    if ( clock_edge == 1'b1 )
    begin: POSEDGE_BLK
      always @(posedge clk)
      begin
        if ( en == enable_active )
        begin
          for (i = 0; i < num_byte_enables; i = i + 1)
          begin
            if ( re[i] == re_active )
              data_out[i*byte_width+: byte_width] <= mem[addr][i*byte_width+: byte_width];
            else
              data_out[i*byte_width+: byte_width] <= {(byte_width){1'bX}};
            if (we[i] == we_active)
              mem[addr][i*byte_width+:byte_width] <= data_in[i*byte_width+:byte_width];
          end
        end
      end
    end else
    begin: NEGEDGE_BLK
      always @(negedge clk)
      begin
        if ( en == enable_active )
        begin
          for (i = 0; i < num_byte_enables; i = i + 1)
          begin
            if ( re[i] == re_active )
              data_out[i*byte_width+: byte_width] <= mem[addr][i*byte_width+: byte_width];
            else
              data_out[i*byte_width+: byte_width] <= {(byte_width){1'bX}};
            if (we[i] == we_active)
              mem[addr][i*byte_width+:byte_width] <= data_in[i*byte_width+:byte_width];
          end
        end
      end
    end
  endgenerate

  // synopsys translate_on

endmodule

module ram_sync_single_be_port ( data_in_d, addr_d, re_d, we_d, data_out_d, data_in, addr, re, we, data_out, clk, a_rst, s_rst, en);

  parameter ram_id = 1;
  parameter words = 16;
  parameter width = 16;
  parameter addr_width = 4;
  parameter [0:0] a_reset_active = 1;
  parameter [0:0] s_reset_active = 1;
  parameter [0:0] enable_active = 1;
  parameter [0:0] re_active = 1;
  parameter [0:0] we_active = 1;
  parameter num_byte_enables = 1;
  parameter [0:0] clock_edge = 1;
  parameter no_of_RAM_readwrite_port = 1;

  input [width-1:0] data_in_d;
  input [addr_width-1:0] addr_d;
  input [num_byte_enables-1:0] re_d;
  input [num_byte_enables-1:0] we_d;
  output [width-1:0] data_out_d;
  output [width-1:0] data_in;
  output [addr_width-1:0] addr;
  output [num_byte_enables-1:0] re;
  output [num_byte_enables-1:0] we;
  input [width-1:0] data_out;
  input clk;
  input a_rst;
  input s_rst;
  input en;

  assign data_in    = data_in_d;
  assign addr       = addr_d;
  assign re         = re_d;
  assign we         = we_d;
  assign data_out_d = data_out;

endmodule

//------> ../td_ccore_solutions/Connections__InBlocking_SysPE__InputType_Connections__SYN_--_e193af7db87ccc7c76c47c5f56a822956142_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:09:55 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  mgc_out_dreg_v2 #(.rscid(32'sd1),
  .width(32'sd8)) data_rsci (
      .d(nl_data_rsci_d[7:0]),
      .z(data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd3),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd329),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__OutBlocking_SysPE__InputType_Connections__SYN--_5dae02d221f0ccc24d0c32e5e6e169c96300_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:09:51 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB_core
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB_core (
  this_val, this_rdy, this_msg, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [7:0] this_msg;
  reg [7:0] this_msg;
  input [7:0] m_rsc_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [7:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire or_dcpl;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  ccs_in_v1 #(.rscid(32'sd4),
  .width(32'sd8)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd6),
  .width(32'sd1)) return_rsci (
      .d(this_rdy),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd328),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  assign or_dcpl = ccs_ccore_start_rsci_idat | asn_itm_1;
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 8'b00000000;
      this_val <= 1'b0;
    end
    else if ( or_dcpl ) begin
      this_msg <= MUX_v_8_2_2(8'b00000000, m_rsci_idat, ccs_ccore_start_rsci_idat);
      this_val <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end

  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB (
  this_val, this_rdy, this_msg, m_rsc_dat, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [7:0] this_msg;
  input [7:0] m_rsc_dat;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB_core Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__InBlocking_SysPE__AccumType_Connections__SYN_--_4a7ec6e3fe4ffbb969ad629169aa89296115_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:09:46 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [31:0] this_msg;
  output [31:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [31:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  mgc_out_dreg_v2 #(.rscid(32'sd7),
  .width(32'sd32)) data_rsci (
      .d(nl_data_rsci_d[31:0]),
      .z(data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd9),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd327),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [31:0] this_msg;
  output [31:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__OutBlocking_SysPE__AccumType_Connections__SYN--_de4c7379377cdb6e2c90db418c7269105beb_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:09:38 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output [31:0] this_msg;
  reg [31:0] this_msg;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire [31:0] m_rsci_idat;
  wire ccs_ccore_start_rsci_idat;
  wire and_dcpl;
  reg io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1;
  wire or_3_cse;
  wire this_val_mx0c1;


  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_ccs_ccore_done_synci_ivld;
  assign nl_ccs_ccore_done_synci_ivld = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1
      & this_rdy;
  ccs_in_v1 #(.rscid(32'sd11),
  .width(32'sd32)) m_rsci (
      .dat(m_rsc_dat),
      .idat(m_rsci_idat)
    );
  ccs_in_v1 #(.rscid(32'sd325),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  ccs_sync_out_vld_v1 #(.rscid(32'sd332)) ccs_ccore_done_synci (
      .vld(ccs_ccore_done_sync_vld),
      .ivld(nl_ccs_ccore_done_synci_ivld[0:0])
    );
  assign or_3_cse = ccs_ccore_start_rsci_idat | and_dcpl;
  assign and_dcpl = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & (~ this_rdy);
  assign this_val_mx0c1 = io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 & this_rdy
      & (~ ccs_ccore_start_rsci_idat);
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( or_3_cse | this_val_mx0c1 ) begin
      this_val <= ~ this_val_mx0c1;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_msg <= 32'b00000000000000000000000000000000;
    end
    else if ( ~(and_dcpl | (~ ccs_ccore_start_rsci_idat)) ) begin
      this_msg <= m_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= 1'b0;
    end
    else begin
      io_read_ccs_ccore_start_rsc_sft_lpi_1_dfm_1 <= or_3_cse;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push
// ------------------------------------------------------------------


module Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push (
  this_val, this_rdy, this_msg, m_rsc_dat, ccs_ccore_start_rsc_dat, ccs_ccore_done_sync_vld,
      ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [31:0] this_msg;
  input [31:0] m_rsc_dat;
  input ccs_ccore_start_rsc_dat;
  output ccs_ccore_done_sync_vld;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .m_rsc_dat(m_rsc_dat),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_ccore_done_sync_vld(ccs_ccore_done_sync_vld),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_SysPE__InputType_Connections__S--_a09193665729a5197eabe9f28a1efa99618f_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:09:34 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB_core
// ------------------------------------------------------------------


module Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB_core
    (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  reg this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  wire [7:0] nl_data_rsci_d;
  assign nl_data_rsci_d = this_msg;
  mgc_out_dreg_v2 #(.rscid(32'sd18),
  .width(32'sd8)) data_rsci (
      .d(nl_data_rsci_d[7:0]),
      .z(data_rsc_z)
    );
  mgc_out_dreg_v2 #(.rscid(32'sd19),
  .width(32'sd1)) return_rsci (
      .d(this_val),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd324),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_rdy <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_rdy <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB
// ------------------------------------------------------------------


module Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB (
  this_val, this_rdy, this_msg, data_rsc_z, return_rsc_z, ccs_ccore_start_rsc_dat,
      ccs_MIO_clk, ccs_MIO_arst
);
  input this_val;
  output this_rdy;
  input [7:0] this_msg;
  output [7:0] data_rsc_z;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB_core Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .this_msg(this_msg),
      .data_rsc_z(data_rsc_z),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
endmodule




//------> ../td_ccore_solutions/Connections__Combinational_SysPE__AccumType_Connections__S--_b0d5d3774c22fe956cb710fa19a5f9a25d23_0/rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:09:30 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB_core
// ------------------------------------------------------------------


module Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB_core
    (
  this_val, this_rdy, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk, ccs_MIO_arst
);
  output this_val;
  reg this_val;
  input this_rdy;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;


  // Interconnect Declarations
  wire ccs_ccore_start_rsci_idat;
  reg asn_itm_1;


  // Interconnect Declarations for Component Instantiations 
  mgc_out_dreg_v2 #(.rscid(32'sd21),
  .width(32'sd1)) return_rsci (
      .d(this_rdy),
      .z(return_rsc_z)
    );
  ccs_in_v1 #(.rscid(32'sd323),
  .width(32'sd1)) ccs_ccore_start_rsci (
      .dat(ccs_ccore_start_rsc_dat),
      .idat(ccs_ccore_start_rsci_idat)
    );
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      this_val <= 1'b0;
    end
    else if ( ccs_ccore_start_rsci_idat | asn_itm_1 ) begin
      this_val <= ccs_ccore_start_rsci_idat;
    end
  end
  always @(posedge ccs_MIO_clk or negedge ccs_MIO_arst) begin
    if ( ~ ccs_MIO_arst ) begin
      asn_itm_1 <= 1'b0;
    end
    else begin
      asn_itm_1 <= ccs_ccore_start_rsci_idat;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB
// ------------------------------------------------------------------


module Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB (
  this_val, this_rdy, this_msg, return_rsc_z, ccs_ccore_start_rsc_dat, ccs_MIO_clk,
      ccs_MIO_arst
);
  output this_val;
  input this_rdy;
  output [31:0] this_msg;
  output return_rsc_z;
  input ccs_ccore_start_rsc_dat;
  input ccs_MIO_clk;
  input ccs_MIO_arst;



  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB_core Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB_core_inst
      (
      .this_val(this_val),
      .this_rdy(this_rdy),
      .return_rsc_z(return_rsc_z),
      .ccs_ccore_start_rsc_dat(ccs_ccore_start_rsc_dat),
      .ccs_MIO_clk(ccs_MIO_clk),
      .ccs_MIO_arst(ccs_MIO_arst)
    );
  assign this_msg = 32'b00000000000000000000000000000000;
endmodule




//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    10.4b/841621 Production Release
//  HLS Date:       Thu Oct 24 17:20:07 PDT 2019
// 
//  Generated by:   billyk@cad.eecs.harvard.edu
//  Generated date: Fri Apr 17 23:29:58 2020
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    SysArray_AccumInRun_AccumInRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysArray_AccumInRun_AccumInRun_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysArray_AccumInRun_AccumInRun_fsm_1
  parameter
    AccumInRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysArray_AccumInRun_AccumInRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // AccumInRun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= AccumInRun_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_ActOutRun_ActOutRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysArray_ActOutRun_ActOutRun_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysArray_ActOutRun_ActOutRun_fsm_1
  parameter
    ActOutRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysArray_ActOutRun_ActOutRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // ActOutRun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= ActOutRun_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_WeightOutRun_WeightOutRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysArray_WeightOutRun_WeightOutRun_fsm (
  clk, rst, fsm_output
);
  input clk;
  input rst;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysArray_WeightOutRun_WeightOutRun_fsm_1
  parameter
    WeightOutRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysArray_WeightOutRun_WeightOutRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // WeightOutRun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= WeightOutRun_rlp_C_0;
    end
    else begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_PERun_fsm
//  FSM Module
// ------------------------------------------------------------------


module SysPE_PERun_PERun_fsm (
  clk, rst, PERun_wen, fsm_output
);
  input clk;
  input rst;
  input PERun_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for SysPE_PERun_PERun_fsm_1
  parameter
    PERun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : SysPE_PERun_PERun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // PERun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= PERun_rlp_C_0;
    end
    else if ( PERun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_staller
// ------------------------------------------------------------------


module SysPE_PERun_staller (
  clk, rst, PERun_wen, PERun_wten, act_out_Push_mioi_wen_comp, accum_out_Push_mioi_wen_comp
);
  input clk;
  input rst;
  output PERun_wen;
  output PERun_wten;
  input act_out_Push_mioi_wen_comp;
  input accum_out_Push_mioi_wen_comp;


  // Interconnect Declarations
  reg PERun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign PERun_wen = act_out_Push_mioi_wen_comp & accum_out_Push_mioi_wen_comp;
  assign PERun_wten = PERun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      PERun_wten_reg <= 1'b0;
    end
    else begin
      PERun_wten_reg <= ~ PERun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp (
  clk, rst, accum_out_Push_mioi_oswt, accum_out_Push_mioi_wen_comp, accum_out_Push_mioi_biwt,
      accum_out_Push_mioi_bdwt, accum_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_wen_comp;
  input accum_out_Push_mioi_biwt;
  input accum_out_Push_mioi_bdwt;
  output accum_out_Push_mioi_bcwt;
  reg accum_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign accum_out_Push_mioi_wen_comp = (~ accum_out_Push_mioi_oswt) | accum_out_Push_mioi_biwt
      | accum_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      accum_out_Push_mioi_bcwt <= ~((~(accum_out_Push_mioi_bcwt | accum_out_Push_mioi_biwt))
          | accum_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl (
  PERun_wen, accum_out_Push_mioi_oswt, accum_out_Push_mioi_biwt, accum_out_Push_mioi_bdwt,
      accum_out_Push_mioi_bcwt, accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct,
      accum_out_Push_mioi_ccs_ccore_done_sync_vld, accum_out_Push_mioi_oswt_pff
);
  input PERun_wen;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_biwt;
  output accum_out_Push_mioi_bdwt;
  input accum_out_Push_mioi_bcwt;
  output accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input accum_out_Push_mioi_ccs_ccore_done_sync_vld;
  input accum_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accum_out_Push_mioi_bdwt = accum_out_Push_mioi_oswt & PERun_wen;
  assign accum_out_Push_mioi_biwt = accum_out_Push_mioi_oswt & (~ accum_out_Push_mioi_bcwt)
      & accum_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct = accum_out_Push_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp (
  clk, rst, act_out_Push_mioi_oswt, act_out_Push_mioi_wen_comp, act_out_Push_mioi_biwt,
      act_out_Push_mioi_bdwt, act_out_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_wen_comp;
  input act_out_Push_mioi_biwt;
  input act_out_Push_mioi_bdwt;
  output act_out_Push_mioi_bcwt;
  reg act_out_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_out_Push_mioi_wen_comp = (~ act_out_Push_mioi_oswt) | act_out_Push_mioi_biwt
      | act_out_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_out_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_out_Push_mioi_bcwt <= ~((~(act_out_Push_mioi_bcwt | act_out_Push_mioi_biwt))
          | act_out_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl (
  PERun_wen, act_out_Push_mioi_oswt, act_out_Push_mioi_biwt, act_out_Push_mioi_bdwt,
      act_out_Push_mioi_bcwt, act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct,
      act_out_Push_mioi_ccs_ccore_done_sync_vld, act_out_Push_mioi_oswt_pff
);
  input PERun_wen;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_biwt;
  output act_out_Push_mioi_bdwt;
  input act_out_Push_mioi_bcwt;
  output act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input act_out_Push_mioi_ccs_ccore_done_sync_vld;
  input act_out_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_out_Push_mioi_bdwt = act_out_Push_mioi_oswt & PERun_wen;
  assign act_out_Push_mioi_biwt = act_out_Push_mioi_oswt & (~ act_out_Push_mioi_bcwt)
      & act_out_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct = act_out_Push_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp (
  clk, rst, accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_in_PopNB_mioi_return_rsc_z_mxwt,
      accum_in_PopNB_mioi_data_rsc_z, accum_in_PopNB_mioi_biwt, accum_in_PopNB_mioi_bdwt,
      accum_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  output accum_in_PopNB_mioi_return_rsc_z_mxwt;
  input [31:0] accum_in_PopNB_mioi_data_rsc_z;
  input accum_in_PopNB_mioi_biwt;
  input accum_in_PopNB_mioi_bdwt;
  input accum_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg accum_in_PopNB_mioi_bcwt;
  reg [31:0] accum_in_PopNB_mioi_data_rsc_z_bfwt;
  reg accum_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign accum_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_32_2_2(accum_in_PopNB_mioi_data_rsc_z,
      accum_in_PopNB_mioi_data_rsc_z_bfwt, accum_in_PopNB_mioi_bcwt);
  assign accum_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(accum_in_PopNB_mioi_return_rsc_z,
      accum_in_PopNB_mioi_return_rsc_z_bfwt, accum_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_in_PopNB_mioi_bcwt <= 1'b0;
      accum_in_PopNB_mioi_data_rsc_z_bfwt <= 32'b00000000000000000000000000000000;
      accum_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      accum_in_PopNB_mioi_bcwt <= ~((~(accum_in_PopNB_mioi_bcwt | accum_in_PopNB_mioi_biwt))
          | accum_in_PopNB_mioi_bdwt);
      accum_in_PopNB_mioi_data_rsc_z_bfwt <= accum_in_PopNB_mioi_data_rsc_z_mxwt;
      accum_in_PopNB_mioi_return_rsc_z_bfwt <= accum_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl (
  PERun_wen, PERun_wten, accum_in_PopNB_mioi_oswt, accum_in_PopNB_mioi_biwt, accum_in_PopNB_mioi_bdwt,
      accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct, accum_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input PERun_wten;
  input accum_in_PopNB_mioi_oswt;
  output accum_in_PopNB_mioi_biwt;
  output accum_in_PopNB_mioi_bdwt;
  output accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input accum_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign accum_in_PopNB_mioi_bdwt = accum_in_PopNB_mioi_oswt & PERun_wen;
  assign accum_in_PopNB_mioi_biwt = (~ PERun_wten) & accum_in_PopNB_mioi_oswt;
  assign accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct = accum_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp (
  clk, rst, act_in_PopNB_mioi_data_rsc_z_mxwt, act_in_PopNB_mioi_return_rsc_z_mxwt,
      act_in_PopNB_mioi_data_rsc_z, act_in_PopNB_mioi_biwt, act_in_PopNB_mioi_bdwt,
      act_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  output act_in_PopNB_mioi_return_rsc_z_mxwt;
  input [7:0] act_in_PopNB_mioi_data_rsc_z;
  input act_in_PopNB_mioi_biwt;
  input act_in_PopNB_mioi_bdwt;
  input act_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg act_in_PopNB_mioi_bcwt;
  reg [7:0] act_in_PopNB_mioi_data_rsc_z_bfwt;
  reg act_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign act_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_8_2_2(act_in_PopNB_mioi_data_rsc_z,
      act_in_PopNB_mioi_data_rsc_z_bfwt, act_in_PopNB_mioi_bcwt);
  assign act_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(act_in_PopNB_mioi_return_rsc_z,
      act_in_PopNB_mioi_return_rsc_z_bfwt, act_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_PopNB_mioi_bcwt <= 1'b0;
      act_in_PopNB_mioi_data_rsc_z_bfwt <= 8'b00000000;
      act_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      act_in_PopNB_mioi_bcwt <= ~((~(act_in_PopNB_mioi_bcwt | act_in_PopNB_mioi_biwt))
          | act_in_PopNB_mioi_bdwt);
      act_in_PopNB_mioi_data_rsc_z_bfwt <= act_in_PopNB_mioi_data_rsc_z_mxwt;
      act_in_PopNB_mioi_return_rsc_z_bfwt <= act_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl (
  PERun_wen, PERun_wten, act_in_PopNB_mioi_oswt, act_in_PopNB_mioi_biwt, act_in_PopNB_mioi_bdwt,
      act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct, act_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input PERun_wten;
  input act_in_PopNB_mioi_oswt;
  output act_in_PopNB_mioi_biwt;
  output act_in_PopNB_mioi_bdwt;
  output act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input act_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_PopNB_mioi_bdwt = act_in_PopNB_mioi_oswt & PERun_wen;
  assign act_in_PopNB_mioi_biwt = (~ PERun_wten) & act_in_PopNB_mioi_oswt;
  assign act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct = act_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_out_PushNB_mioi_weight_out_PushNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_weight_out_PushNB_mioi_weight_out_PushNB_mio_wait_ctrl (
  PERun_wten, weight_out_PushNB_mioi_iswt0, weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct
);
  input PERun_wten;
  input weight_out_PushNB_mioi_iswt0;
  output weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;



  // Interconnect Declarations for Component Instantiations 
  assign weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct = weight_out_PushNB_mioi_iswt0
      & (~ PERun_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp (
  clk, rst, weight_in_PopNB_mioi_data_rsc_z_mxwt, weight_in_PopNB_mioi_return_rsc_z_mxwt,
      weight_in_PopNB_mioi_data_rsc_z, weight_in_PopNB_mioi_biwt, weight_in_PopNB_mioi_bdwt,
      weight_in_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  output weight_in_PopNB_mioi_return_rsc_z_mxwt;
  input [7:0] weight_in_PopNB_mioi_data_rsc_z;
  input weight_in_PopNB_mioi_biwt;
  input weight_in_PopNB_mioi_bdwt;
  input weight_in_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg weight_in_PopNB_mioi_bcwt;
  reg [7:0] weight_in_PopNB_mioi_data_rsc_z_bfwt;
  reg weight_in_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign weight_in_PopNB_mioi_data_rsc_z_mxwt = MUX_v_8_2_2(weight_in_PopNB_mioi_data_rsc_z,
      weight_in_PopNB_mioi_data_rsc_z_bfwt, weight_in_PopNB_mioi_bcwt);
  assign weight_in_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(weight_in_PopNB_mioi_return_rsc_z,
      weight_in_PopNB_mioi_return_rsc_z_bfwt, weight_in_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_in_PopNB_mioi_bcwt <= 1'b0;
      weight_in_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      weight_in_PopNB_mioi_bcwt <= ~((~(weight_in_PopNB_mioi_bcwt | weight_in_PopNB_mioi_biwt))
          | weight_in_PopNB_mioi_bdwt);
      weight_in_PopNB_mioi_return_rsc_z_bfwt <= weight_in_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_in_PopNB_mioi_data_rsc_z_bfwt <= 8'b00000000;
    end
    else if ( ~ weight_in_PopNB_mioi_bcwt ) begin
      weight_in_PopNB_mioi_data_rsc_z_bfwt <= weight_in_PopNB_mioi_data_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl (
  PERun_wen, weight_in_PopNB_mioi_oswt, PERun_wten, weight_in_PopNB_mioi_biwt, weight_in_PopNB_mioi_bdwt,
      weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct, weight_in_PopNB_mioi_oswt_pff
);
  input PERun_wen;
  input weight_in_PopNB_mioi_oswt;
  input PERun_wten;
  output weight_in_PopNB_mioi_biwt;
  output weight_in_PopNB_mioi_bdwt;
  output weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  input weight_in_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign weight_in_PopNB_mioi_bdwt = weight_in_PopNB_mioi_oswt & PERun_wen;
  assign weight_in_PopNB_mioi_biwt = (~ PERun_wten) & weight_in_PopNB_mioi_oswt;
  assign weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct = weight_in_PopNB_mioi_oswt_pff
      & PERun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_304_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
// ------------------------------------------------------------------


module InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_304_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
    (
  en, data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d,
      en_d
);
  output en;
  input [7:0] data_out;
  output we;
  output re;
  output [4:0] addr;
  output [7:0] data_in;
  input [7:0] data_in_d;
  input [4:0] addr_d;
  input re_d;
  input we_d;
  output [7:0] data_out_d;
  input en_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_303_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
// ------------------------------------------------------------------


module InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_303_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
    (
  en, data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d,
      en_d
);
  output en;
  input [7:0] data_out;
  output we;
  output re;
  output [4:0] addr;
  output [7:0] data_in;
  input [7:0] data_in_d;
  input [4:0] addr_d;
  input re_d;
  input we_d;
  output [7:0] data_out_d;
  input en_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_302_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
// ------------------------------------------------------------------


module InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_302_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
    (
  en, data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d,
      en_d
);
  output en;
  input [7:0] data_out;
  output we;
  output re;
  output [4:0] addr;
  output [7:0] data_in;
  input [7:0] data_in_d;
  input [4:0] addr_d;
  input re_d;
  input we_d;
  output [7:0] data_out_d;
  input en_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_301_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
// ------------------------------------------------------------------


module InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_301_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
    (
  en, data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d,
      en_d
);
  output en;
  input [7:0] data_out;
  output we;
  output re;
  output [4:0] addr;
  output [7:0] data_in;
  input [7:0] data_in_d;
  input [4:0] addr_d;
  input re_d;
  input we_d;
  output [7:0] data_out_d;
  input en_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_300_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
// ------------------------------------------------------------------


module InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_300_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
    (
  en, data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d,
      en_d
);
  output en;
  input [7:0] data_out;
  output we;
  output re;
  output [4:0] addr;
  output [7:0] data_in;
  input [7:0] data_in_d;
  input [4:0] addr_d;
  input re_d;
  input we_d;
  output [7:0] data_out_d;
  input en_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_299_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
// ------------------------------------------------------------------


module InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_299_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
    (
  en, data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d,
      en_d
);
  output en;
  input [7:0] data_out;
  output we;
  output re;
  output [4:0] addr;
  output [7:0] data_in;
  input [7:0] data_in_d;
  input [4:0] addr_d;
  input re_d;
  input we_d;
  output [7:0] data_out_d;
  input en_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_298_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
// ------------------------------------------------------------------


module InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_298_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
    (
  en, data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d,
      en_d
);
  output en;
  input [7:0] data_out;
  output we;
  output re;
  output [4:0] addr;
  output [7:0] data_in;
  input [7:0] data_in_d;
  input [4:0] addr_d;
  input re_d;
  input we_d;
  output [7:0] data_out_d;
  input en_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_297_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
// ------------------------------------------------------------------


module InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_297_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
    (
  en, data_out, we, re, addr, data_in, data_in_d, addr_d, re_d, we_d, data_out_d,
      en_d
);
  output en;
  input [7:0] data_out;
  output we;
  output re;
  output [4:0] addr;
  output [7:0] data_in;
  input [7:0] data_in_d;
  input [4:0] addr_d;
  input re_d;
  input we_d;
  output [7:0] data_out_d;
  input en_d;



  // Interconnect Declarations for Component Instantiations 
  assign en = (en_d);
  assign data_out_d = data_out;
  assign we = (we_d);
  assign re = (re_d);
  assign addr = (addr_d);
  assign data_in = (data_in_d);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_ReadRspRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_ReadRspRun_fsm (
  clk, rst, ReadRspRun_wen, fsm_output
);
  input clk;
  input rst;
  input ReadRspRun_wen;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for InputSetup_ReadRspRun_ReadRspRun_fsm_1
  parameter
    ReadRspRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputSetup_ReadRspRun_ReadRspRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // ReadRspRun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= ReadRspRun_rlp_C_0;
    end
    else if ( ReadRspRun_wen ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_staller_2
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_staller_2 (
  clk, rst, ReadRspRun_wen, ReadRspRun_wten, act_in_vec_Push_mioi_wen_comp, act_in_vec_Push_1_mioi_wen_comp,
      act_in_vec_Push_2_mioi_wen_comp, act_in_vec_Push_3_mioi_wen_comp, act_in_vec_Push_4_mioi_wen_comp,
      act_in_vec_Push_5_mioi_wen_comp, act_in_vec_Push_6_mioi_wen_comp, act_in_vec_Push_7_mioi_wen_comp
);
  input clk;
  input rst;
  output ReadRspRun_wen;
  output ReadRspRun_wten;
  input act_in_vec_Push_mioi_wen_comp;
  input act_in_vec_Push_1_mioi_wen_comp;
  input act_in_vec_Push_2_mioi_wen_comp;
  input act_in_vec_Push_3_mioi_wen_comp;
  input act_in_vec_Push_4_mioi_wen_comp;
  input act_in_vec_Push_5_mioi_wen_comp;
  input act_in_vec_Push_6_mioi_wen_comp;
  input act_in_vec_Push_7_mioi_wen_comp;


  // Interconnect Declarations
  reg ReadRspRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign ReadRspRun_wen = act_in_vec_Push_mioi_wen_comp & act_in_vec_Push_1_mioi_wen_comp
      & act_in_vec_Push_2_mioi_wen_comp & act_in_vec_Push_3_mioi_wen_comp & act_in_vec_Push_4_mioi_wen_comp
      & act_in_vec_Push_5_mioi_wen_comp & act_in_vec_Push_6_mioi_wen_comp & act_in_vec_Push_7_mioi_wen_comp;
  assign ReadRspRun_wten = ReadRspRun_wten_reg;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      ReadRspRun_wten_reg <= 1'b0;
    end
    else begin
      ReadRspRun_wten_reg <= ~ ReadRspRun_wen;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_act_in_vec_Push_7_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_act_in_vec_Push_7_mio_wait_dp
    (
  clk, rst, act_in_vec_Push_7_mioi_oswt, act_in_vec_Push_7_mioi_wen_comp, act_in_vec_Push_7_mioi_biwt,
      act_in_vec_Push_7_mioi_bdwt, act_in_vec_Push_7_mioi_bcwt
);
  input clk;
  input rst;
  input act_in_vec_Push_7_mioi_oswt;
  output act_in_vec_Push_7_mioi_wen_comp;
  input act_in_vec_Push_7_mioi_biwt;
  input act_in_vec_Push_7_mioi_bdwt;
  output act_in_vec_Push_7_mioi_bcwt;
  reg act_in_vec_Push_7_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_7_mioi_wen_comp = (~ act_in_vec_Push_7_mioi_oswt) | act_in_vec_Push_7_mioi_biwt
      | act_in_vec_Push_7_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_vec_Push_7_mioi_bcwt <= 1'b0;
    end
    else begin
      act_in_vec_Push_7_mioi_bcwt <= ~((~(act_in_vec_Push_7_mioi_bcwt | act_in_vec_Push_7_mioi_biwt))
          | act_in_vec_Push_7_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_act_in_vec_Push_7_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_act_in_vec_Push_7_mio_wait_ctrl
    (
  ReadRspRun_wen, act_in_vec_Push_7_mioi_oswt, act_in_vec_Push_7_mioi_biwt, act_in_vec_Push_7_mioi_bdwt,
      act_in_vec_Push_7_mioi_bcwt, act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      act_in_vec_Push_7_mioi_ccs_ccore_done_sync_vld, act_in_vec_Push_7_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input act_in_vec_Push_7_mioi_oswt;
  output act_in_vec_Push_7_mioi_biwt;
  output act_in_vec_Push_7_mioi_bdwt;
  input act_in_vec_Push_7_mioi_bcwt;
  output act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input act_in_vec_Push_7_mioi_ccs_ccore_done_sync_vld;
  input act_in_vec_Push_7_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_7_mioi_bdwt = act_in_vec_Push_7_mioi_oswt & ReadRspRun_wen;
  assign act_in_vec_Push_7_mioi_biwt = act_in_vec_Push_7_mioi_oswt & (~ act_in_vec_Push_7_mioi_bcwt)
      & act_in_vec_Push_7_mioi_ccs_ccore_done_sync_vld;
  assign act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = act_in_vec_Push_7_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_act_in_vec_Push_6_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_act_in_vec_Push_6_mio_wait_dp
    (
  clk, rst, act_in_vec_Push_6_mioi_oswt, act_in_vec_Push_6_mioi_wen_comp, act_in_vec_Push_6_mioi_biwt,
      act_in_vec_Push_6_mioi_bdwt, act_in_vec_Push_6_mioi_bcwt
);
  input clk;
  input rst;
  input act_in_vec_Push_6_mioi_oswt;
  output act_in_vec_Push_6_mioi_wen_comp;
  input act_in_vec_Push_6_mioi_biwt;
  input act_in_vec_Push_6_mioi_bdwt;
  output act_in_vec_Push_6_mioi_bcwt;
  reg act_in_vec_Push_6_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_6_mioi_wen_comp = (~ act_in_vec_Push_6_mioi_oswt) | act_in_vec_Push_6_mioi_biwt
      | act_in_vec_Push_6_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_vec_Push_6_mioi_bcwt <= 1'b0;
    end
    else begin
      act_in_vec_Push_6_mioi_bcwt <= ~((~(act_in_vec_Push_6_mioi_bcwt | act_in_vec_Push_6_mioi_biwt))
          | act_in_vec_Push_6_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_act_in_vec_Push_6_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_act_in_vec_Push_6_mio_wait_ctrl
    (
  ReadRspRun_wen, act_in_vec_Push_6_mioi_oswt, act_in_vec_Push_6_mioi_biwt, act_in_vec_Push_6_mioi_bdwt,
      act_in_vec_Push_6_mioi_bcwt, act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      act_in_vec_Push_6_mioi_ccs_ccore_done_sync_vld, act_in_vec_Push_6_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input act_in_vec_Push_6_mioi_oswt;
  output act_in_vec_Push_6_mioi_biwt;
  output act_in_vec_Push_6_mioi_bdwt;
  input act_in_vec_Push_6_mioi_bcwt;
  output act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input act_in_vec_Push_6_mioi_ccs_ccore_done_sync_vld;
  input act_in_vec_Push_6_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_6_mioi_bdwt = act_in_vec_Push_6_mioi_oswt & ReadRspRun_wen;
  assign act_in_vec_Push_6_mioi_biwt = act_in_vec_Push_6_mioi_oswt & (~ act_in_vec_Push_6_mioi_bcwt)
      & act_in_vec_Push_6_mioi_ccs_ccore_done_sync_vld;
  assign act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = act_in_vec_Push_6_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_act_in_vec_Push_5_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_act_in_vec_Push_5_mio_wait_dp
    (
  clk, rst, act_in_vec_Push_5_mioi_oswt, act_in_vec_Push_5_mioi_wen_comp, act_in_vec_Push_5_mioi_biwt,
      act_in_vec_Push_5_mioi_bdwt, act_in_vec_Push_5_mioi_bcwt
);
  input clk;
  input rst;
  input act_in_vec_Push_5_mioi_oswt;
  output act_in_vec_Push_5_mioi_wen_comp;
  input act_in_vec_Push_5_mioi_biwt;
  input act_in_vec_Push_5_mioi_bdwt;
  output act_in_vec_Push_5_mioi_bcwt;
  reg act_in_vec_Push_5_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_5_mioi_wen_comp = (~ act_in_vec_Push_5_mioi_oswt) | act_in_vec_Push_5_mioi_biwt
      | act_in_vec_Push_5_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_vec_Push_5_mioi_bcwt <= 1'b0;
    end
    else begin
      act_in_vec_Push_5_mioi_bcwt <= ~((~(act_in_vec_Push_5_mioi_bcwt | act_in_vec_Push_5_mioi_biwt))
          | act_in_vec_Push_5_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_act_in_vec_Push_5_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_act_in_vec_Push_5_mio_wait_ctrl
    (
  ReadRspRun_wen, act_in_vec_Push_5_mioi_oswt, act_in_vec_Push_5_mioi_biwt, act_in_vec_Push_5_mioi_bdwt,
      act_in_vec_Push_5_mioi_bcwt, act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      act_in_vec_Push_5_mioi_ccs_ccore_done_sync_vld, act_in_vec_Push_5_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input act_in_vec_Push_5_mioi_oswt;
  output act_in_vec_Push_5_mioi_biwt;
  output act_in_vec_Push_5_mioi_bdwt;
  input act_in_vec_Push_5_mioi_bcwt;
  output act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input act_in_vec_Push_5_mioi_ccs_ccore_done_sync_vld;
  input act_in_vec_Push_5_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_5_mioi_bdwt = act_in_vec_Push_5_mioi_oswt & ReadRspRun_wen;
  assign act_in_vec_Push_5_mioi_biwt = act_in_vec_Push_5_mioi_oswt & (~ act_in_vec_Push_5_mioi_bcwt)
      & act_in_vec_Push_5_mioi_ccs_ccore_done_sync_vld;
  assign act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = act_in_vec_Push_5_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_act_in_vec_Push_4_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_act_in_vec_Push_4_mio_wait_dp
    (
  clk, rst, act_in_vec_Push_4_mioi_oswt, act_in_vec_Push_4_mioi_wen_comp, act_in_vec_Push_4_mioi_biwt,
      act_in_vec_Push_4_mioi_bdwt, act_in_vec_Push_4_mioi_bcwt
);
  input clk;
  input rst;
  input act_in_vec_Push_4_mioi_oswt;
  output act_in_vec_Push_4_mioi_wen_comp;
  input act_in_vec_Push_4_mioi_biwt;
  input act_in_vec_Push_4_mioi_bdwt;
  output act_in_vec_Push_4_mioi_bcwt;
  reg act_in_vec_Push_4_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_4_mioi_wen_comp = (~ act_in_vec_Push_4_mioi_oswt) | act_in_vec_Push_4_mioi_biwt
      | act_in_vec_Push_4_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_vec_Push_4_mioi_bcwt <= 1'b0;
    end
    else begin
      act_in_vec_Push_4_mioi_bcwt <= ~((~(act_in_vec_Push_4_mioi_bcwt | act_in_vec_Push_4_mioi_biwt))
          | act_in_vec_Push_4_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_act_in_vec_Push_4_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_act_in_vec_Push_4_mio_wait_ctrl
    (
  ReadRspRun_wen, act_in_vec_Push_4_mioi_oswt, act_in_vec_Push_4_mioi_biwt, act_in_vec_Push_4_mioi_bdwt,
      act_in_vec_Push_4_mioi_bcwt, act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      act_in_vec_Push_4_mioi_ccs_ccore_done_sync_vld, act_in_vec_Push_4_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input act_in_vec_Push_4_mioi_oswt;
  output act_in_vec_Push_4_mioi_biwt;
  output act_in_vec_Push_4_mioi_bdwt;
  input act_in_vec_Push_4_mioi_bcwt;
  output act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input act_in_vec_Push_4_mioi_ccs_ccore_done_sync_vld;
  input act_in_vec_Push_4_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_4_mioi_bdwt = act_in_vec_Push_4_mioi_oswt & ReadRspRun_wen;
  assign act_in_vec_Push_4_mioi_biwt = act_in_vec_Push_4_mioi_oswt & (~ act_in_vec_Push_4_mioi_bcwt)
      & act_in_vec_Push_4_mioi_ccs_ccore_done_sync_vld;
  assign act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = act_in_vec_Push_4_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_act_in_vec_Push_3_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_act_in_vec_Push_3_mio_wait_dp
    (
  clk, rst, act_in_vec_Push_3_mioi_oswt, act_in_vec_Push_3_mioi_wen_comp, act_in_vec_Push_3_mioi_biwt,
      act_in_vec_Push_3_mioi_bdwt, act_in_vec_Push_3_mioi_bcwt
);
  input clk;
  input rst;
  input act_in_vec_Push_3_mioi_oswt;
  output act_in_vec_Push_3_mioi_wen_comp;
  input act_in_vec_Push_3_mioi_biwt;
  input act_in_vec_Push_3_mioi_bdwt;
  output act_in_vec_Push_3_mioi_bcwt;
  reg act_in_vec_Push_3_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_3_mioi_wen_comp = (~ act_in_vec_Push_3_mioi_oswt) | act_in_vec_Push_3_mioi_biwt
      | act_in_vec_Push_3_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_vec_Push_3_mioi_bcwt <= 1'b0;
    end
    else begin
      act_in_vec_Push_3_mioi_bcwt <= ~((~(act_in_vec_Push_3_mioi_bcwt | act_in_vec_Push_3_mioi_biwt))
          | act_in_vec_Push_3_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_act_in_vec_Push_3_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_act_in_vec_Push_3_mio_wait_ctrl
    (
  ReadRspRun_wen, act_in_vec_Push_3_mioi_oswt, act_in_vec_Push_3_mioi_biwt, act_in_vec_Push_3_mioi_bdwt,
      act_in_vec_Push_3_mioi_bcwt, act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      act_in_vec_Push_3_mioi_ccs_ccore_done_sync_vld, act_in_vec_Push_3_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input act_in_vec_Push_3_mioi_oswt;
  output act_in_vec_Push_3_mioi_biwt;
  output act_in_vec_Push_3_mioi_bdwt;
  input act_in_vec_Push_3_mioi_bcwt;
  output act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input act_in_vec_Push_3_mioi_ccs_ccore_done_sync_vld;
  input act_in_vec_Push_3_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_3_mioi_bdwt = act_in_vec_Push_3_mioi_oswt & ReadRspRun_wen;
  assign act_in_vec_Push_3_mioi_biwt = act_in_vec_Push_3_mioi_oswt & (~ act_in_vec_Push_3_mioi_bcwt)
      & act_in_vec_Push_3_mioi_ccs_ccore_done_sync_vld;
  assign act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = act_in_vec_Push_3_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_act_in_vec_Push_2_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_act_in_vec_Push_2_mio_wait_dp
    (
  clk, rst, act_in_vec_Push_2_mioi_oswt, act_in_vec_Push_2_mioi_wen_comp, act_in_vec_Push_2_mioi_biwt,
      act_in_vec_Push_2_mioi_bdwt, act_in_vec_Push_2_mioi_bcwt
);
  input clk;
  input rst;
  input act_in_vec_Push_2_mioi_oswt;
  output act_in_vec_Push_2_mioi_wen_comp;
  input act_in_vec_Push_2_mioi_biwt;
  input act_in_vec_Push_2_mioi_bdwt;
  output act_in_vec_Push_2_mioi_bcwt;
  reg act_in_vec_Push_2_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_2_mioi_wen_comp = (~ act_in_vec_Push_2_mioi_oswt) | act_in_vec_Push_2_mioi_biwt
      | act_in_vec_Push_2_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_vec_Push_2_mioi_bcwt <= 1'b0;
    end
    else begin
      act_in_vec_Push_2_mioi_bcwt <= ~((~(act_in_vec_Push_2_mioi_bcwt | act_in_vec_Push_2_mioi_biwt))
          | act_in_vec_Push_2_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_act_in_vec_Push_2_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_act_in_vec_Push_2_mio_wait_ctrl
    (
  ReadRspRun_wen, act_in_vec_Push_2_mioi_oswt, act_in_vec_Push_2_mioi_biwt, act_in_vec_Push_2_mioi_bdwt,
      act_in_vec_Push_2_mioi_bcwt, act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      act_in_vec_Push_2_mioi_ccs_ccore_done_sync_vld, act_in_vec_Push_2_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input act_in_vec_Push_2_mioi_oswt;
  output act_in_vec_Push_2_mioi_biwt;
  output act_in_vec_Push_2_mioi_bdwt;
  input act_in_vec_Push_2_mioi_bcwt;
  output act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input act_in_vec_Push_2_mioi_ccs_ccore_done_sync_vld;
  input act_in_vec_Push_2_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_2_mioi_bdwt = act_in_vec_Push_2_mioi_oswt & ReadRspRun_wen;
  assign act_in_vec_Push_2_mioi_biwt = act_in_vec_Push_2_mioi_oswt & (~ act_in_vec_Push_2_mioi_bcwt)
      & act_in_vec_Push_2_mioi_ccs_ccore_done_sync_vld;
  assign act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = act_in_vec_Push_2_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_act_in_vec_Push_1_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_act_in_vec_Push_1_mio_wait_dp
    (
  clk, rst, act_in_vec_Push_1_mioi_oswt, act_in_vec_Push_1_mioi_wen_comp, act_in_vec_Push_1_mioi_biwt,
      act_in_vec_Push_1_mioi_bdwt, act_in_vec_Push_1_mioi_bcwt
);
  input clk;
  input rst;
  input act_in_vec_Push_1_mioi_oswt;
  output act_in_vec_Push_1_mioi_wen_comp;
  input act_in_vec_Push_1_mioi_biwt;
  input act_in_vec_Push_1_mioi_bdwt;
  output act_in_vec_Push_1_mioi_bcwt;
  reg act_in_vec_Push_1_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_1_mioi_wen_comp = (~ act_in_vec_Push_1_mioi_oswt) | act_in_vec_Push_1_mioi_biwt
      | act_in_vec_Push_1_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_vec_Push_1_mioi_bcwt <= 1'b0;
    end
    else begin
      act_in_vec_Push_1_mioi_bcwt <= ~((~(act_in_vec_Push_1_mioi_bcwt | act_in_vec_Push_1_mioi_biwt))
          | act_in_vec_Push_1_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_act_in_vec_Push_1_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_act_in_vec_Push_1_mio_wait_ctrl
    (
  ReadRspRun_wen, act_in_vec_Push_1_mioi_oswt, act_in_vec_Push_1_mioi_biwt, act_in_vec_Push_1_mioi_bdwt,
      act_in_vec_Push_1_mioi_bcwt, act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      act_in_vec_Push_1_mioi_ccs_ccore_done_sync_vld, act_in_vec_Push_1_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input act_in_vec_Push_1_mioi_oswt;
  output act_in_vec_Push_1_mioi_biwt;
  output act_in_vec_Push_1_mioi_bdwt;
  input act_in_vec_Push_1_mioi_bcwt;
  output act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input act_in_vec_Push_1_mioi_ccs_ccore_done_sync_vld;
  input act_in_vec_Push_1_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_1_mioi_bdwt = act_in_vec_Push_1_mioi_oswt & ReadRspRun_wen;
  assign act_in_vec_Push_1_mioi_biwt = act_in_vec_Push_1_mioi_oswt & (~ act_in_vec_Push_1_mioi_bcwt)
      & act_in_vec_Push_1_mioi_ccs_ccore_done_sync_vld;
  assign act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = act_in_vec_Push_1_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_mioi_act_in_vec_Push_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_mioi_act_in_vec_Push_mio_wait_dp (
  clk, rst, act_in_vec_Push_mioi_oswt, act_in_vec_Push_mioi_wen_comp, act_in_vec_Push_mioi_biwt,
      act_in_vec_Push_mioi_bdwt, act_in_vec_Push_mioi_bcwt
);
  input clk;
  input rst;
  input act_in_vec_Push_mioi_oswt;
  output act_in_vec_Push_mioi_wen_comp;
  input act_in_vec_Push_mioi_biwt;
  input act_in_vec_Push_mioi_bdwt;
  output act_in_vec_Push_mioi_bcwt;
  reg act_in_vec_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_mioi_wen_comp = (~ act_in_vec_Push_mioi_oswt) | act_in_vec_Push_mioi_biwt
      | act_in_vec_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_in_vec_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      act_in_vec_Push_mioi_bcwt <= ~((~(act_in_vec_Push_mioi_bcwt | act_in_vec_Push_mioi_biwt))
          | act_in_vec_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_mioi_act_in_vec_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_mioi_act_in_vec_Push_mio_wait_ctrl (
  ReadRspRun_wen, act_in_vec_Push_mioi_oswt, act_in_vec_Push_mioi_biwt, act_in_vec_Push_mioi_bdwt,
      act_in_vec_Push_mioi_bcwt, act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      act_in_vec_Push_mioi_ccs_ccore_done_sync_vld, act_in_vec_Push_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input act_in_vec_Push_mioi_oswt;
  output act_in_vec_Push_mioi_biwt;
  output act_in_vec_Push_mioi_bdwt;
  input act_in_vec_Push_mioi_bcwt;
  output act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input act_in_vec_Push_mioi_ccs_ccore_done_sync_vld;
  input act_in_vec_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign act_in_vec_Push_mioi_bdwt = act_in_vec_Push_mioi_oswt & ReadRspRun_wen;
  assign act_in_vec_Push_mioi_biwt = act_in_vec_Push_mioi_oswt & (~ act_in_vec_Push_mioi_bcwt)
      & act_in_vec_Push_mioi_ccs_ccore_done_sync_vld;
  assign act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = act_in_vec_Push_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_rsp_inter_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_rsp_inter_PopNB_mio_wait_dp (
  clk, rst, rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt, rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt,
      rsp_inter_PopNB_mioi_return_rsc_z_mxwt, rsp_inter_PopNB_mioi_data_valids_rsc_z,
      rsp_inter_PopNB_mioi_biwt, rsp_inter_PopNB_mioi_bdwt, rsp_inter_PopNB_mioi_data_data_rsc_z,
      rsp_inter_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [7:0] rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
  output [63:0] rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt;
  output rsp_inter_PopNB_mioi_return_rsc_z_mxwt;
  input [7:0] rsp_inter_PopNB_mioi_data_valids_rsc_z;
  input rsp_inter_PopNB_mioi_biwt;
  input rsp_inter_PopNB_mioi_bdwt;
  input [63:0] rsp_inter_PopNB_mioi_data_data_rsc_z;
  input rsp_inter_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg rsp_inter_PopNB_mioi_bcwt;
  reg [7:0] rsp_inter_PopNB_mioi_data_valids_rsc_z_bfwt;
  reg [63:0] rsp_inter_PopNB_mioi_data_data_rsc_z_bfwt;
  reg rsp_inter_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt = MUX_v_8_2_2(rsp_inter_PopNB_mioi_data_valids_rsc_z,
      rsp_inter_PopNB_mioi_data_valids_rsc_z_bfwt, rsp_inter_PopNB_mioi_bcwt);
  assign rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_64_2_2(rsp_inter_PopNB_mioi_data_data_rsc_z,
      rsp_inter_PopNB_mioi_data_data_rsc_z_bfwt, rsp_inter_PopNB_mioi_bcwt);
  assign rsp_inter_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(rsp_inter_PopNB_mioi_return_rsc_z,
      rsp_inter_PopNB_mioi_return_rsc_z_bfwt, rsp_inter_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rsp_inter_PopNB_mioi_bcwt <= 1'b0;
      rsp_inter_PopNB_mioi_data_valids_rsc_z_bfwt <= 8'b00000000;
      rsp_inter_PopNB_mioi_data_data_rsc_z_bfwt <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      rsp_inter_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      rsp_inter_PopNB_mioi_bcwt <= ~((~(rsp_inter_PopNB_mioi_bcwt | rsp_inter_PopNB_mioi_biwt))
          | rsp_inter_PopNB_mioi_bdwt);
      rsp_inter_PopNB_mioi_data_valids_rsc_z_bfwt <= rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
      rsp_inter_PopNB_mioi_data_data_rsc_z_bfwt <= rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt;
      rsp_inter_PopNB_mioi_return_rsc_z_bfwt <= rsp_inter_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_rsp_inter_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_rsp_inter_PopNB_mio_wait_ctrl (
  ReadRspRun_wen, rsp_inter_PopNB_mioi_oswt, ReadRspRun_wten, rsp_inter_PopNB_mioi_biwt,
      rsp_inter_PopNB_mioi_bdwt, rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct,
      rsp_inter_PopNB_mioi_oswt_pff
);
  input ReadRspRun_wen;
  input rsp_inter_PopNB_mioi_oswt;
  input ReadRspRun_wten;
  output rsp_inter_PopNB_mioi_biwt;
  output rsp_inter_PopNB_mioi_bdwt;
  output rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  input rsp_inter_PopNB_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rsp_inter_PopNB_mioi_bdwt = rsp_inter_PopNB_mioi_oswt & ReadRspRun_wen;
  assign rsp_inter_PopNB_mioi_biwt = (~ ReadRspRun_wten) & rsp_inter_PopNB_mioi_oswt;
  assign rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct = rsp_inter_PopNB_mioi_oswt_pff
      & ReadRspRun_wen;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadReqRun_ReadReqRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputSetup_ReadReqRun_ReadReqRun_fsm (
  clk, rst, start_Pop_mioi_wen_comp, fsm_output, while_C_1_tr0, while_if_for_C_1_tr0
);
  input clk;
  input rst;
  input start_Pop_mioi_wen_comp;
  output [5:0] fsm_output;
  reg [5:0] fsm_output;
  input while_C_1_tr0;
  input while_if_for_C_1_tr0;


  // FSM State Type Declaration for InputSetup_ReadReqRun_ReadReqRun_fsm_1
  parameter
    ReadReqRun_rlp_C_0 = 3'd0,
    while_C_0 = 3'd1,
    while_C_1 = 3'd2,
    while_if_for_C_0 = 3'd3,
    while_if_for_C_1 = 3'd4,
    while_C_2 = 3'd5;

  reg [2:0] state_var;
  reg [2:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputSetup_ReadReqRun_ReadReqRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 6'b000010;
        state_var_NS = while_C_1;
      end
      while_C_1 : begin
        fsm_output = 6'b000100;
        if ( while_C_1_tr0 ) begin
          state_var_NS = while_C_2;
        end
        else begin
          state_var_NS = while_if_for_C_0;
        end
      end
      while_if_for_C_0 : begin
        fsm_output = 6'b001000;
        state_var_NS = while_if_for_C_1;
      end
      while_if_for_C_1 : begin
        fsm_output = 6'b010000;
        if ( while_if_for_C_1_tr0 ) begin
          state_var_NS = while_C_2;
        end
        else begin
          state_var_NS = while_if_for_C_0;
        end
      end
      while_C_2 : begin
        fsm_output = 6'b100000;
        state_var_NS = while_C_0;
      end
      // ReadReqRun_rlp_C_0
      default : begin
        fsm_output = 6'b000001;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= ReadReqRun_rlp_C_0;
    end
    else if ( start_Pop_mioi_wen_comp ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadReqRun_staller_1
// ------------------------------------------------------------------


module InputSetup_ReadReqRun_staller_1 (
  start_Pop_mioi_wen_comp, ReadReqRun_wten_pff
);
  input start_Pop_mioi_wen_comp;
  output ReadReqRun_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign ReadReqRun_wten_pff = ~ start_Pop_mioi_wen_comp;
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadReqRun_req_inter_PushNB_mioi_req_inter_PushNB_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadReqRun_req_inter_PushNB_mioi_req_inter_PushNB_mio_wait_ctrl
    (
  req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_pff, req_inter_PushNB_mioi_iswt0_pff,
      ReadReqRun_wten_pff
);
  output req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_pff;
  input req_inter_PushNB_mioi_iswt0_pff;
  input ReadReqRun_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_pff = req_inter_PushNB_mioi_iswt0_pff
      & (~ ReadReqRun_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadReqRun_start_Pop_mioi_start_Pop_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_ReadReqRun_start_Pop_mioi_start_Pop_mio_wait_dp (
  clk, rst, start_Pop_mioi_oswt, start_Pop_mioi_wen_comp, start_Pop_mioi_biwt, start_Pop_mioi_bdwt,
      start_Pop_mioi_bcwt
);
  input clk;
  input rst;
  input start_Pop_mioi_oswt;
  output start_Pop_mioi_wen_comp;
  input start_Pop_mioi_biwt;
  input start_Pop_mioi_bdwt;
  output start_Pop_mioi_bcwt;
  reg start_Pop_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign start_Pop_mioi_wen_comp = (~ start_Pop_mioi_oswt) | start_Pop_mioi_biwt
      | start_Pop_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      start_Pop_mioi_bcwt <= 1'b0;
    end
    else begin
      start_Pop_mioi_bcwt <= ~((~(start_Pop_mioi_bcwt | start_Pop_mioi_biwt)) | start_Pop_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadReqRun_start_Pop_mioi_start_Pop_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_ReadReqRun_start_Pop_mioi_start_Pop_mio_wait_ctrl (
  ReadReqRun_wen, start_Pop_mioi_oswt, ReadReqRun_wten, start_Pop_mioi_biwt, start_Pop_mioi_bdwt,
      start_Pop_mioi_bcwt, start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_sct,
      start_Pop_mioi_ccs_ccore_done_sync_vld, start_Pop_mioi_oswt_pff
);
  input ReadReqRun_wen;
  input start_Pop_mioi_oswt;
  input ReadReqRun_wten;
  output start_Pop_mioi_biwt;
  output start_Pop_mioi_bdwt;
  input start_Pop_mioi_bcwt;
  output start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_sct;
  input start_Pop_mioi_ccs_ccore_done_sync_vld;
  input start_Pop_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign start_Pop_mioi_bdwt = start_Pop_mioi_oswt & ReadReqRun_wen;
  assign start_Pop_mioi_biwt = start_Pop_mioi_oswt & (~ start_Pop_mioi_bcwt) & start_Pop_mioi_ccs_ccore_done_sync_vld;
  assign start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_sct = start_Pop_mioi_oswt_pff
      & (~ ReadReqRun_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_MemoryRun_fsm
//  FSM Module
// ------------------------------------------------------------------


module InputSetup_MemoryRun_MemoryRun_fsm (
  clk, rst, rsp_inter_Push_mioi_wen_comp, fsm_output
);
  input clk;
  input rst;
  input rsp_inter_Push_mioi_wen_comp;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;


  // FSM State Type Declaration for InputSetup_MemoryRun_MemoryRun_fsm_1
  parameter
    MemoryRun_rlp_C_0 = 1'd0,
    while_C_0 = 1'd1;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : InputSetup_MemoryRun_MemoryRun_fsm_1
    case (state_var)
      while_C_0 : begin
        fsm_output = 2'b10;
        state_var_NS = while_C_0;
      end
      // MemoryRun_rlp_C_0
      default : begin
        fsm_output = 2'b01;
        state_var_NS = while_C_0;
      end
    endcase
  end

  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      state_var <= MemoryRun_rlp_C_0;
    end
    else if ( rsp_inter_Push_mioi_wen_comp ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_staller
// ------------------------------------------------------------------


module InputSetup_MemoryRun_staller (
  clk, rst, MemoryRun_wten, rsp_inter_Push_mioi_wen_comp, MemoryRun_wten_pff
);
  input clk;
  input rst;
  output MemoryRun_wten;
  input rsp_inter_Push_mioi_wen_comp;
  output MemoryRun_wten_pff;


  // Interconnect Declarations
  reg MemoryRun_wten_reg;


  // Interconnect Declarations for Component Instantiations 
  assign MemoryRun_wten = MemoryRun_wten_reg;
  assign MemoryRun_wten_pff = ~ rsp_inter_Push_mioi_wen_comp;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      MemoryRun_wten_reg <= 1'b0;
    end
    else begin
      MemoryRun_wten_reg <= ~ rsp_inter_Push_mioi_wen_comp;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_wait_dp
// ------------------------------------------------------------------


module InputSetup_MemoryRun_wait_dp (
  clk, rst, mem_inst_banks_bank_array_impl_data0_rsc_cgo_iro, mem_inst_banks_bank_array_impl_data0_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data0_rsci_en_d, mem_inst_banks_bank_array_impl_data1_rsc_cgo_iro,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d, mem_inst_banks_bank_array_impl_data1_rsci_en_d,
      mem_inst_banks_bank_array_impl_data2_rsc_cgo_iro, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data2_rsci_en_d, mem_inst_banks_bank_array_impl_data3_rsc_cgo_iro,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d, mem_inst_banks_bank_array_impl_data3_rsci_en_d,
      mem_inst_banks_bank_array_impl_data4_rsc_cgo_iro, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data4_rsci_en_d, mem_inst_banks_bank_array_impl_data5_rsc_cgo_iro,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d, mem_inst_banks_bank_array_impl_data5_rsci_en_d,
      mem_inst_banks_bank_array_impl_data6_rsc_cgo_iro, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data6_rsci_en_d, mem_inst_banks_bank_array_impl_data7_rsc_cgo_iro,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d, mem_inst_banks_bank_array_impl_data7_rsci_en_d,
      MemoryRun_wen, mem_inst_banks_bank_array_impl_data0_rsc_cgo, mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsc_cgo, mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data2_rsc_cgo, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsc_cgo, mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data4_rsc_cgo, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsc_cgo, mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data6_rsc_cgo, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsc_cgo, mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg
);
  input clk;
  input rst;
  input mem_inst_banks_bank_array_impl_data0_rsc_cgo_iro;
  input [7:0] mem_inst_banks_bank_array_impl_data0_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data0_rsci_en_d;
  input mem_inst_banks_bank_array_impl_data1_rsc_cgo_iro;
  input [7:0] mem_inst_banks_bank_array_impl_data1_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data1_rsci_en_d;
  input mem_inst_banks_bank_array_impl_data2_rsc_cgo_iro;
  input [7:0] mem_inst_banks_bank_array_impl_data2_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data2_rsci_en_d;
  input mem_inst_banks_bank_array_impl_data3_rsc_cgo_iro;
  input [7:0] mem_inst_banks_bank_array_impl_data3_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data3_rsci_en_d;
  input mem_inst_banks_bank_array_impl_data4_rsc_cgo_iro;
  input [7:0] mem_inst_banks_bank_array_impl_data4_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data4_rsci_en_d;
  input mem_inst_banks_bank_array_impl_data5_rsc_cgo_iro;
  input [7:0] mem_inst_banks_bank_array_impl_data5_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data5_rsci_en_d;
  input mem_inst_banks_bank_array_impl_data6_rsc_cgo_iro;
  input [7:0] mem_inst_banks_bank_array_impl_data6_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data6_rsci_en_d;
  input mem_inst_banks_bank_array_impl_data7_rsc_cgo_iro;
  input [7:0] mem_inst_banks_bank_array_impl_data7_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data7_rsci_en_d;
  input MemoryRun_wen;
  input mem_inst_banks_bank_array_impl_data0_rsc_cgo;
  output [7:0] mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg;
  reg [7:0] mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg;
  input mem_inst_banks_bank_array_impl_data1_rsc_cgo;
  output [7:0] mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg;
  reg [7:0] mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg;
  input mem_inst_banks_bank_array_impl_data2_rsc_cgo;
  output [7:0] mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg;
  reg [7:0] mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg;
  input mem_inst_banks_bank_array_impl_data3_rsc_cgo;
  output [7:0] mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg;
  reg [7:0] mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg;
  input mem_inst_banks_bank_array_impl_data4_rsc_cgo;
  output [7:0] mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg;
  reg [7:0] mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg;
  input mem_inst_banks_bank_array_impl_data5_rsc_cgo;
  output [7:0] mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg;
  reg [7:0] mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg;
  input mem_inst_banks_bank_array_impl_data6_rsc_cgo;
  output [7:0] mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg;
  reg [7:0] mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg;
  input mem_inst_banks_bank_array_impl_data7_rsc_cgo;
  output [7:0] mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg;
  reg [7:0] mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg;



  // Interconnect Declarations for Component Instantiations 
  assign mem_inst_banks_bank_array_impl_data0_rsci_en_d = ~(MemoryRun_wen & (mem_inst_banks_bank_array_impl_data0_rsc_cgo
      | mem_inst_banks_bank_array_impl_data0_rsc_cgo_iro));
  assign mem_inst_banks_bank_array_impl_data1_rsci_en_d = ~(MemoryRun_wen & (mem_inst_banks_bank_array_impl_data1_rsc_cgo
      | mem_inst_banks_bank_array_impl_data1_rsc_cgo_iro));
  assign mem_inst_banks_bank_array_impl_data2_rsci_en_d = ~(MemoryRun_wen & (mem_inst_banks_bank_array_impl_data2_rsc_cgo
      | mem_inst_banks_bank_array_impl_data2_rsc_cgo_iro));
  assign mem_inst_banks_bank_array_impl_data3_rsci_en_d = ~(MemoryRun_wen & (mem_inst_banks_bank_array_impl_data3_rsc_cgo
      | mem_inst_banks_bank_array_impl_data3_rsc_cgo_iro));
  assign mem_inst_banks_bank_array_impl_data4_rsci_en_d = ~(MemoryRun_wen & (mem_inst_banks_bank_array_impl_data4_rsc_cgo
      | mem_inst_banks_bank_array_impl_data4_rsc_cgo_iro));
  assign mem_inst_banks_bank_array_impl_data5_rsci_en_d = ~(MemoryRun_wen & (mem_inst_banks_bank_array_impl_data5_rsc_cgo
      | mem_inst_banks_bank_array_impl_data5_rsc_cgo_iro));
  assign mem_inst_banks_bank_array_impl_data6_rsci_en_d = ~(MemoryRun_wen & (mem_inst_banks_bank_array_impl_data6_rsc_cgo
      | mem_inst_banks_bank_array_impl_data6_rsc_cgo_iro));
  assign mem_inst_banks_bank_array_impl_data7_rsci_en_d = ~(MemoryRun_wen & (mem_inst_banks_bank_array_impl_data7_rsc_cgo
      | mem_inst_banks_bank_array_impl_data7_rsc_cgo_iro));
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg <= 8'b00000000;
    end
    else if ( ~ mem_inst_banks_bank_array_impl_data0_rsci_en_d ) begin
      mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg <= mem_inst_banks_bank_array_impl_data0_rsci_data_out_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg <= 8'b00000000;
    end
    else if ( ~ mem_inst_banks_bank_array_impl_data1_rsci_en_d ) begin
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg <= mem_inst_banks_bank_array_impl_data1_rsci_data_out_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg <= 8'b00000000;
    end
    else if ( ~ mem_inst_banks_bank_array_impl_data2_rsci_en_d ) begin
      mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg <= mem_inst_banks_bank_array_impl_data2_rsci_data_out_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg <= 8'b00000000;
    end
    else if ( ~ mem_inst_banks_bank_array_impl_data3_rsci_en_d ) begin
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg <= mem_inst_banks_bank_array_impl_data3_rsci_data_out_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg <= 8'b00000000;
    end
    else if ( ~ mem_inst_banks_bank_array_impl_data4_rsci_en_d ) begin
      mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg <= mem_inst_banks_bank_array_impl_data4_rsci_data_out_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg <= 8'b00000000;
    end
    else if ( ~ mem_inst_banks_bank_array_impl_data5_rsci_en_d ) begin
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg <= mem_inst_banks_bank_array_impl_data5_rsci_data_out_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg <= 8'b00000000;
    end
    else if ( ~ mem_inst_banks_bank_array_impl_data6_rsci_en_d ) begin
      mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg <= mem_inst_banks_bank_array_impl_data6_rsci_data_out_d;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg <= 8'b00000000;
    end
    else if ( ~ mem_inst_banks_bank_array_impl_data7_rsci_en_d ) begin
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg <= mem_inst_banks_bank_array_impl_data7_rsci_data_out_d;
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_rsp_inter_Push_mioi_rsp_inter_Push_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_MemoryRun_rsp_inter_Push_mioi_rsp_inter_Push_mio_wait_dp (
  clk, rst, rsp_inter_Push_mioi_oswt, rsp_inter_Push_mioi_wen_comp, rsp_inter_Push_mioi_biwt,
      rsp_inter_Push_mioi_bdwt, rsp_inter_Push_mioi_bcwt
);
  input clk;
  input rst;
  input rsp_inter_Push_mioi_oswt;
  output rsp_inter_Push_mioi_wen_comp;
  input rsp_inter_Push_mioi_biwt;
  input rsp_inter_Push_mioi_bdwt;
  output rsp_inter_Push_mioi_bcwt;
  reg rsp_inter_Push_mioi_bcwt;



  // Interconnect Declarations for Component Instantiations 
  assign rsp_inter_Push_mioi_wen_comp = (~ rsp_inter_Push_mioi_oswt) | rsp_inter_Push_mioi_biwt
      | rsp_inter_Push_mioi_bcwt;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      rsp_inter_Push_mioi_bcwt <= 1'b0;
    end
    else begin
      rsp_inter_Push_mioi_bcwt <= ~((~(rsp_inter_Push_mioi_bcwt | rsp_inter_Push_mioi_biwt))
          | rsp_inter_Push_mioi_bdwt);
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_rsp_inter_Push_mioi_rsp_inter_Push_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_MemoryRun_rsp_inter_Push_mioi_rsp_inter_Push_mio_wait_ctrl (
  MemoryRun_wen, MemoryRun_wten, rsp_inter_Push_mioi_oswt, rsp_inter_Push_mioi_biwt,
      rsp_inter_Push_mioi_bdwt, rsp_inter_Push_mioi_bcwt, rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct,
      rsp_inter_Push_mioi_ccs_ccore_done_sync_vld, rsp_inter_Push_mioi_oswt_pff
);
  input MemoryRun_wen;
  input MemoryRun_wten;
  input rsp_inter_Push_mioi_oswt;
  output rsp_inter_Push_mioi_biwt;
  output rsp_inter_Push_mioi_bdwt;
  input rsp_inter_Push_mioi_bcwt;
  output rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct;
  input rsp_inter_Push_mioi_ccs_ccore_done_sync_vld;
  input rsp_inter_Push_mioi_oswt_pff;



  // Interconnect Declarations for Component Instantiations 
  assign rsp_inter_Push_mioi_bdwt = rsp_inter_Push_mioi_oswt & MemoryRun_wen;
  assign rsp_inter_Push_mioi_biwt = rsp_inter_Push_mioi_oswt & (~ rsp_inter_Push_mioi_bcwt)
      & rsp_inter_Push_mioi_ccs_ccore_done_sync_vld;
  assign rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct = rsp_inter_Push_mioi_oswt_pff
      & (~ MemoryRun_wten);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_write_req_PopNB_mioi_write_req_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_MemoryRun_write_req_PopNB_mioi_write_req_PopNB_mio_wait_dp (
  clk, rst, write_req_PopNB_mioi_data_data_data_rsc_z_mxwt, write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      write_req_PopNB_mioi_return_rsc_z_mxwt, write_req_PopNB_mioi_data_data_data_rsc_z,
      write_req_PopNB_mioi_biwt, write_req_PopNB_mioi_bdwt, write_req_PopNB_mioi_data_index_rsc_z,
      write_req_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output [63:0] write_req_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [4:0] write_req_PopNB_mioi_data_index_rsc_z_mxwt;
  output write_req_PopNB_mioi_return_rsc_z_mxwt;
  input [63:0] write_req_PopNB_mioi_data_data_data_rsc_z;
  input write_req_PopNB_mioi_biwt;
  input write_req_PopNB_mioi_bdwt;
  input [4:0] write_req_PopNB_mioi_data_index_rsc_z;
  input write_req_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg write_req_PopNB_mioi_bcwt;
  reg [63:0] write_req_PopNB_mioi_data_data_data_rsc_z_bfwt;
  reg [4:0] write_req_PopNB_mioi_data_index_rsc_z_bfwt;
  reg write_req_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign write_req_PopNB_mioi_data_data_data_rsc_z_mxwt = MUX_v_64_2_2(write_req_PopNB_mioi_data_data_data_rsc_z,
      write_req_PopNB_mioi_data_data_data_rsc_z_bfwt, write_req_PopNB_mioi_bcwt);
  assign write_req_PopNB_mioi_data_index_rsc_z_mxwt = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z,
      write_req_PopNB_mioi_data_index_rsc_z_bfwt, write_req_PopNB_mioi_bcwt);
  assign write_req_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(write_req_PopNB_mioi_return_rsc_z,
      write_req_PopNB_mioi_return_rsc_z_bfwt, write_req_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      write_req_PopNB_mioi_bcwt <= 1'b0;
      write_req_PopNB_mioi_data_data_data_rsc_z_bfwt <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      write_req_PopNB_mioi_data_index_rsc_z_bfwt <= 5'b00000;
      write_req_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      write_req_PopNB_mioi_bcwt <= ~((~(write_req_PopNB_mioi_bcwt | write_req_PopNB_mioi_biwt))
          | write_req_PopNB_mioi_bdwt);
      write_req_PopNB_mioi_data_data_data_rsc_z_bfwt <= write_req_PopNB_mioi_data_data_data_rsc_z_mxwt;
      write_req_PopNB_mioi_data_index_rsc_z_bfwt <= write_req_PopNB_mioi_data_index_rsc_z_mxwt;
      write_req_PopNB_mioi_return_rsc_z_bfwt <= write_req_PopNB_mioi_return_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_write_req_PopNB_mioi_write_req_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_MemoryRun_write_req_PopNB_mioi_write_req_PopNB_mio_wait_ctrl (
  MemoryRun_wen, MemoryRun_wten, write_req_PopNB_mioi_oswt, write_req_PopNB_mioi_biwt,
      write_req_PopNB_mioi_bdwt, write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct,
      write_req_PopNB_mioi_oswt_pff, MemoryRun_wten_pff
);
  input MemoryRun_wen;
  input MemoryRun_wten;
  input write_req_PopNB_mioi_oswt;
  output write_req_PopNB_mioi_biwt;
  output write_req_PopNB_mioi_bdwt;
  output write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct;
  input write_req_PopNB_mioi_oswt_pff;
  input MemoryRun_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign write_req_PopNB_mioi_bdwt = write_req_PopNB_mioi_oswt & MemoryRun_wen;
  assign write_req_PopNB_mioi_biwt = (~ MemoryRun_wten) & write_req_PopNB_mioi_oswt;
  assign write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct = write_req_PopNB_mioi_oswt_pff
      & (~ MemoryRun_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_req_inter_PopNB_mioi_req_inter_PopNB_mio_wait_dp
// ------------------------------------------------------------------


module InputSetup_MemoryRun_req_inter_PopNB_mioi_req_inter_PopNB_mio_wait_dp (
  clk, rst, req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt, req_inter_PopNB_mioi_data_valids_rsc_z_mxwt,
      req_inter_PopNB_mioi_data_addr_rsc_z_mxwt, req_inter_PopNB_mioi_data_data_rsc_z_mxwt,
      req_inter_PopNB_mioi_return_rsc_z_mxwt, req_inter_PopNB_mioi_data_type_val_rsc_z,
      req_inter_PopNB_mioi_biwt, req_inter_PopNB_mioi_bdwt, req_inter_PopNB_mioi_data_valids_rsc_z,
      req_inter_PopNB_mioi_data_addr_rsc_z, req_inter_PopNB_mioi_data_data_rsc_z,
      req_inter_PopNB_mioi_return_rsc_z
);
  input clk;
  input rst;
  output req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt;
  output [7:0] req_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
  output [63:0] req_inter_PopNB_mioi_data_addr_rsc_z_mxwt;
  output [63:0] req_inter_PopNB_mioi_data_data_rsc_z_mxwt;
  output req_inter_PopNB_mioi_return_rsc_z_mxwt;
  input req_inter_PopNB_mioi_data_type_val_rsc_z;
  input req_inter_PopNB_mioi_biwt;
  input req_inter_PopNB_mioi_bdwt;
  input [7:0] req_inter_PopNB_mioi_data_valids_rsc_z;
  input [63:0] req_inter_PopNB_mioi_data_addr_rsc_z;
  input [63:0] req_inter_PopNB_mioi_data_data_rsc_z;
  input req_inter_PopNB_mioi_return_rsc_z;


  // Interconnect Declarations
  reg req_inter_PopNB_mioi_bcwt;
  reg req_inter_PopNB_mioi_data_type_val_rsc_z_bfwt;
  reg [7:0] req_inter_PopNB_mioi_data_valids_rsc_z_bfwt;
  reg [63:0] req_inter_PopNB_mioi_data_addr_rsc_z_bfwt;
  reg [63:0] req_inter_PopNB_mioi_data_data_rsc_z_bfwt;
  reg req_inter_PopNB_mioi_return_rsc_z_bfwt;


  // Interconnect Declarations for Component Instantiations 
  assign req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt = MUX_s_1_2_2(req_inter_PopNB_mioi_data_type_val_rsc_z,
      req_inter_PopNB_mioi_data_type_val_rsc_z_bfwt, req_inter_PopNB_mioi_bcwt);
  assign req_inter_PopNB_mioi_data_valids_rsc_z_mxwt = MUX_v_8_2_2(req_inter_PopNB_mioi_data_valids_rsc_z,
      req_inter_PopNB_mioi_data_valids_rsc_z_bfwt, req_inter_PopNB_mioi_bcwt);
  assign req_inter_PopNB_mioi_data_addr_rsc_z_mxwt = MUX_v_64_2_2(req_inter_PopNB_mioi_data_addr_rsc_z,
      req_inter_PopNB_mioi_data_addr_rsc_z_bfwt, req_inter_PopNB_mioi_bcwt);
  assign req_inter_PopNB_mioi_data_data_rsc_z_mxwt = MUX_v_64_2_2(req_inter_PopNB_mioi_data_data_rsc_z,
      req_inter_PopNB_mioi_data_data_rsc_z_bfwt, req_inter_PopNB_mioi_bcwt);
  assign req_inter_PopNB_mioi_return_rsc_z_mxwt = MUX_s_1_2_2(req_inter_PopNB_mioi_return_rsc_z,
      req_inter_PopNB_mioi_return_rsc_z_bfwt, req_inter_PopNB_mioi_bcwt);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      req_inter_PopNB_mioi_bcwt <= 1'b0;
      req_inter_PopNB_mioi_data_type_val_rsc_z_bfwt <= 1'b0;
      req_inter_PopNB_mioi_return_rsc_z_bfwt <= 1'b0;
    end
    else begin
      req_inter_PopNB_mioi_bcwt <= ~((~(req_inter_PopNB_mioi_bcwt | req_inter_PopNB_mioi_biwt))
          | req_inter_PopNB_mioi_bdwt);
      req_inter_PopNB_mioi_data_type_val_rsc_z_bfwt <= req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt;
      req_inter_PopNB_mioi_return_rsc_z_bfwt <= req_inter_PopNB_mioi_return_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      req_inter_PopNB_mioi_data_valids_rsc_z_bfwt <= 8'b00000000;
    end
    else if ( ~ req_inter_PopNB_mioi_bcwt ) begin
      req_inter_PopNB_mioi_data_valids_rsc_z_bfwt <= req_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      req_inter_PopNB_mioi_data_addr_rsc_z_bfwt <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ req_inter_PopNB_mioi_bcwt ) begin
      req_inter_PopNB_mioi_data_addr_rsc_z_bfwt <= req_inter_PopNB_mioi_data_addr_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      req_inter_PopNB_mioi_data_data_rsc_z_bfwt <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
    end
    else if ( ~ req_inter_PopNB_mioi_bcwt ) begin
      req_inter_PopNB_mioi_data_data_rsc_z_bfwt <= req_inter_PopNB_mioi_data_data_rsc_z_mxwt;
    end
  end

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [63:0] MUX_v_64_2_2;
    input [63:0] input_0;
    input [63:0] input_1;
    input [0:0] sel;
    reg [63:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_64_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_req_inter_PopNB_mioi_req_inter_PopNB_mio_wait_ctrl
// ------------------------------------------------------------------


module InputSetup_MemoryRun_req_inter_PopNB_mioi_req_inter_PopNB_mio_wait_ctrl (
  MemoryRun_wen, req_inter_PopNB_mioi_oswt, MemoryRun_wten, req_inter_PopNB_mioi_biwt,
      req_inter_PopNB_mioi_bdwt, req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct,
      req_inter_PopNB_mioi_oswt_pff, MemoryRun_wten_pff
);
  input MemoryRun_wen;
  input req_inter_PopNB_mioi_oswt;
  input MemoryRun_wten;
  output req_inter_PopNB_mioi_biwt;
  output req_inter_PopNB_mioi_bdwt;
  output req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct;
  input req_inter_PopNB_mioi_oswt_pff;
  input MemoryRun_wten_pff;



  // Interconnect Declarations for Component Instantiations 
  assign req_inter_PopNB_mioi_bdwt = req_inter_PopNB_mioi_oswt & MemoryRun_wen;
  assign req_inter_PopNB_mioi_biwt = (~ MemoryRun_wten) & req_inter_PopNB_mioi_oswt;
  assign req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct = req_inter_PopNB_mioi_oswt_pff
      & (~ MemoryRun_wten_pff);
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_AccumInRun
// ------------------------------------------------------------------


module SysArray_AccumInRun (
  clk, rst, accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_pff
);
  input clk;
  input rst;
  output accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_pff;


  // Interconnect Declarations
  wire [1:0] fsm_output;

  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_1;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_2;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_3;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_4;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_5;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_6;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_7;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7;

  // Interconnect Declarations for Component Instantiations 
  SysArray_AccumInRun_AccumInRun_fsm SysArray_AccumInRun_AccumInRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign p0_Unreachable_virtual_function_in_abstract_class_prb = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb  -> p0_Unreachable_virtual_function_in_abstract_class_prb );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_1 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_1 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1  -> p0_Unreachable_virtual_function_in_abstract_class_prb_1 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_2 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_2 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2  -> p0_Unreachable_virtual_function_in_abstract_class_prb_2 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_3 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_3 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3  -> p0_Unreachable_virtual_function_in_abstract_class_prb_3 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_4 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_4 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4  -> p0_Unreachable_virtual_function_in_abstract_class_prb_4 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_5 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_5 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5  -> p0_Unreachable_virtual_function_in_abstract_class_prb_5 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_6 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_6 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6  -> p0_Unreachable_virtual_function_in_abstract_class_prb_6 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_7 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 3314
  // psl default clock = (posedge clk);
  // psl SysArray_AccumInRun_connections_h_ln3314_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_7 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7  -> p0_Unreachable_virtual_function_in_abstract_class_prb_7 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7 = 1'b0;
  assign accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_pff = fsm_output[1];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_ActOutRun
// ------------------------------------------------------------------


module SysArray_ActOutRun (
  clk, rst, act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_pff
);
  input clk;
  input rst;
  output act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_pff;


  // Interconnect Declarations
  wire [1:0] fsm_output;


  // Interconnect Declarations for Component Instantiations 
  SysArray_ActOutRun_ActOutRun_fsm SysArray_ActOutRun_ActOutRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_pff = fsm_output[1];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray_WeightOutRun
// ------------------------------------------------------------------


module SysArray_WeightOutRun (
  clk, rst, weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_pff
);
  input clk;
  input rst;
  output weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_pff;


  // Interconnect Declarations
  wire [1:0] fsm_output;


  // Interconnect Declarations for Component Instantiations 
  SysArray_WeightOutRun_WeightOutRun_fsm SysArray_WeightOutRun_WeightOutRun_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .fsm_output(fsm_output)
    );
  assign weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_pff = fsm_output[1];
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_out_Push_mioi
// ------------------------------------------------------------------


module SysPE_PERun_accum_out_Push_mioi (
  clk, rst, accum_out_val, accum_out_rdy, accum_out_msg, PERun_wen, accum_out_Push_mioi_oswt,
      accum_out_Push_mioi_wen_comp, accum_out_Push_mioi_m_rsc_dat_PERun, accum_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;
  input PERun_wen;
  input accum_out_Push_mioi_oswt;
  output accum_out_Push_mioi_wen_comp;
  input [31:0] accum_out_Push_mioi_m_rsc_dat_PERun;
  input accum_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire accum_out_Push_mioi_biwt;
  wire accum_out_Push_mioi_bdwt;
  wire accum_out_Push_mioi_bcwt;
  wire accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  wire accum_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_AccumType_Connections_SYN_PORT_Push  accum_out_Push_mioi
      (
      .this_val(accum_out_val),
      .this_rdy(accum_out_rdy),
      .this_msg(accum_out_msg),
      .m_rsc_dat(accum_out_Push_mioi_m_rsc_dat_PERun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .ccs_ccore_done_sync_vld(accum_out_Push_mioi_ccs_ccore_done_sync_vld)
    );
  SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .accum_out_Push_mioi_oswt(accum_out_Push_mioi_oswt),
      .accum_out_Push_mioi_biwt(accum_out_Push_mioi_biwt),
      .accum_out_Push_mioi_bdwt(accum_out_Push_mioi_bdwt),
      .accum_out_Push_mioi_bcwt(accum_out_Push_mioi_bcwt),
      .accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct(accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .accum_out_Push_mioi_ccs_ccore_done_sync_vld(accum_out_Push_mioi_ccs_ccore_done_sync_vld),
      .accum_out_Push_mioi_oswt_pff(accum_out_Push_mioi_oswt_pff)
    );
  SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp SysPE_PERun_accum_out_Push_mioi_accum_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .accum_out_Push_mioi_oswt(accum_out_Push_mioi_oswt),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_biwt(accum_out_Push_mioi_biwt),
      .accum_out_Push_mioi_bdwt(accum_out_Push_mioi_bdwt),
      .accum_out_Push_mioi_bcwt(accum_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_out_Push_mioi
// ------------------------------------------------------------------


module SysPE_PERun_act_out_Push_mioi (
  clk, rst, act_out_val, act_out_rdy, act_out_msg, PERun_wen, act_out_Push_mioi_oswt,
      act_out_Push_mioi_wen_comp, act_out_Push_mioi_m_rsc_dat_PERun, act_out_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  input PERun_wen;
  input act_out_Push_mioi_oswt;
  output act_out_Push_mioi_wen_comp;
  input [7:0] act_out_Push_mioi_m_rsc_dat_PERun;
  input act_out_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_out_Push_mioi_biwt;
  wire act_out_Push_mioi_bdwt;
  wire act_out_Push_mioi_bcwt;
  wire act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct;
  wire act_out_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_out_Push_mioi
      (
      .this_val(act_out_val),
      .this_rdy(act_out_rdy),
      .this_msg(act_out_msg),
      .m_rsc_dat(act_out_Push_mioi_m_rsc_dat_PERun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .ccs_ccore_done_sync_vld(act_out_Push_mioi_ccs_ccore_done_sync_vld)
    );
  SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .act_out_Push_mioi_oswt(act_out_Push_mioi_oswt),
      .act_out_Push_mioi_biwt(act_out_Push_mioi_biwt),
      .act_out_Push_mioi_bdwt(act_out_Push_mioi_bdwt),
      .act_out_Push_mioi_bcwt(act_out_Push_mioi_bcwt),
      .act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct(act_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .act_out_Push_mioi_ccs_ccore_done_sync_vld(act_out_Push_mioi_ccs_ccore_done_sync_vld),
      .act_out_Push_mioi_oswt_pff(act_out_Push_mioi_oswt_pff)
    );
  SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp SysPE_PERun_act_out_Push_mioi_act_out_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_out_Push_mioi_oswt(act_out_Push_mioi_oswt),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .act_out_Push_mioi_biwt(act_out_Push_mioi_biwt),
      .act_out_Push_mioi_bdwt(act_out_Push_mioi_bdwt),
      .act_out_Push_mioi_bcwt(act_out_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_accum_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_accum_in_PopNB_mioi (
  clk, rst, accum_in_val, accum_in_rdy, accum_in_msg, PERun_wen, PERun_wten, accum_in_PopNB_mioi_oswt,
      accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_in_PopNB_mioi_return_rsc_z_mxwt,
      accum_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  input PERun_wen;
  input PERun_wten;
  input accum_in_PopNB_mioi_oswt;
  output [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  output accum_in_PopNB_mioi_return_rsc_z_mxwt;
  input accum_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [31:0] accum_in_PopNB_mioi_data_rsc_z;
  wire accum_in_PopNB_mioi_biwt;
  wire accum_in_PopNB_mioi_bdwt;
  wire accum_in_PopNB_mioi_return_rsc_z;
  wire accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_AccumType_Connections_SYN_PORT_PopNB  accum_in_PopNB_mioi
      (
      .this_val(accum_in_val),
      .this_rdy(accum_in_rdy),
      .this_msg(accum_in_msg),
      .data_rsc_z(accum_in_PopNB_mioi_data_rsc_z),
      .return_rsc_z(accum_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
  SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .accum_in_PopNB_mioi_oswt(accum_in_PopNB_mioi_oswt),
      .accum_in_PopNB_mioi_biwt(accum_in_PopNB_mioi_biwt),
      .accum_in_PopNB_mioi_bdwt(accum_in_PopNB_mioi_bdwt),
      .accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct(accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .accum_in_PopNB_mioi_oswt_pff(accum_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp SysPE_PERun_accum_in_PopNB_mioi_accum_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .accum_in_PopNB_mioi_data_rsc_z_mxwt(accum_in_PopNB_mioi_data_rsc_z_mxwt),
      .accum_in_PopNB_mioi_return_rsc_z_mxwt(accum_in_PopNB_mioi_return_rsc_z_mxwt),
      .accum_in_PopNB_mioi_data_rsc_z(accum_in_PopNB_mioi_data_rsc_z),
      .accum_in_PopNB_mioi_biwt(accum_in_PopNB_mioi_biwt),
      .accum_in_PopNB_mioi_bdwt(accum_in_PopNB_mioi_bdwt),
      .accum_in_PopNB_mioi_return_rsc_z(accum_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_act_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_act_in_PopNB_mioi (
  clk, rst, act_in_val, act_in_rdy, act_in_msg, PERun_wen, PERun_wten, act_in_PopNB_mioi_oswt,
      act_in_PopNB_mioi_data_rsc_z_mxwt, act_in_PopNB_mioi_return_rsc_z_mxwt, act_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input PERun_wen;
  input PERun_wten;
  input act_in_PopNB_mioi_oswt;
  output [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  output act_in_PopNB_mioi_return_rsc_z_mxwt;
  input act_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [7:0] act_in_PopNB_mioi_data_rsc_z;
  wire act_in_PopNB_mioi_biwt;
  wire act_in_PopNB_mioi_bdwt;
  wire act_in_PopNB_mioi_return_rsc_z;
  wire act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB  act_in_PopNB_mioi
      (
      .this_val(act_in_val),
      .this_rdy(act_in_rdy),
      .this_msg(act_in_msg),
      .data_rsc_z(act_in_PopNB_mioi_data_rsc_z),
      .return_rsc_z(act_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
  SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_in_PopNB_mioi_oswt(act_in_PopNB_mioi_oswt),
      .act_in_PopNB_mioi_biwt(act_in_PopNB_mioi_biwt),
      .act_in_PopNB_mioi_bdwt(act_in_PopNB_mioi_bdwt),
      .act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct(act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .act_in_PopNB_mioi_oswt_pff(act_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp SysPE_PERun_act_in_PopNB_mioi_act_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_PopNB_mioi_data_rsc_z_mxwt(act_in_PopNB_mioi_data_rsc_z_mxwt),
      .act_in_PopNB_mioi_return_rsc_z_mxwt(act_in_PopNB_mioi_return_rsc_z_mxwt),
      .act_in_PopNB_mioi_data_rsc_z(act_in_PopNB_mioi_data_rsc_z),
      .act_in_PopNB_mioi_biwt(act_in_PopNB_mioi_biwt),
      .act_in_PopNB_mioi_bdwt(act_in_PopNB_mioi_bdwt),
      .act_in_PopNB_mioi_return_rsc_z(act_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_out_PushNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_weight_out_PushNB_mioi (
  clk, rst, weight_out_val, weight_out_rdy, weight_out_msg, PERun_wten, weight_out_PushNB_mioi_iswt0,
      weight_out_PushNB_mioi_m_rsc_dat_PERun
);
  input clk;
  input rst;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;
  input PERun_wten;
  input weight_out_PushNB_mioi_iswt0;
  input [7:0] weight_out_PushNB_mioi_m_rsc_dat_PERun;


  // Interconnect Declarations
  wire weight_out_PushNB_mioi_return_rsc_z;
  wire weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_PushNB  weight_out_PushNB_mioi
      (
      .this_val(weight_out_val),
      .this_rdy(weight_out_rdy),
      .this_msg(weight_out_msg),
      .m_rsc_dat(weight_out_PushNB_mioi_m_rsc_dat_PERun),
      .return_rsc_z(weight_out_PushNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
  SysPE_PERun_weight_out_PushNB_mioi_weight_out_PushNB_mio_wait_ctrl SysPE_PERun_weight_out_PushNB_mioi_weight_out_PushNB_mio_wait_ctrl_inst
      (
      .PERun_wten(PERun_wten),
      .weight_out_PushNB_mioi_iswt0(weight_out_PushNB_mioi_iswt0),
      .weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct(weight_out_PushNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun_weight_in_PopNB_mioi
// ------------------------------------------------------------------


module SysPE_PERun_weight_in_PopNB_mioi (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, PERun_wen, weight_in_PopNB_mioi_oswt,
      PERun_wten, weight_in_PopNB_mioi_data_rsc_z_mxwt, weight_in_PopNB_mioi_return_rsc_z_mxwt,
      weight_in_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input PERun_wen;
  input weight_in_PopNB_mioi_oswt;
  input PERun_wten;
  output [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  output weight_in_PopNB_mioi_return_rsc_z_mxwt;
  input weight_in_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [7:0] weight_in_PopNB_mioi_data_rsc_z;
  wire weight_in_PopNB_mioi_biwt;
  wire weight_in_PopNB_mioi_bdwt;
  wire weight_in_PopNB_mioi_return_rsc_z;
  wire weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_in_PopNB_mioi
      (
      .this_val(weight_in_val),
      .this_rdy(weight_in_rdy),
      .this_msg(weight_in_msg),
      .data_rsc_z(weight_in_PopNB_mioi_data_rsc_z),
      .return_rsc_z(weight_in_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct)
    );
  SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_ctrl_inst
      (
      .PERun_wen(PERun_wen),
      .weight_in_PopNB_mioi_oswt(weight_in_PopNB_mioi_oswt),
      .PERun_wten(PERun_wten),
      .weight_in_PopNB_mioi_biwt(weight_in_PopNB_mioi_biwt),
      .weight_in_PopNB_mioi_bdwt(weight_in_PopNB_mioi_bdwt),
      .weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct(weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_sct),
      .weight_in_PopNB_mioi_oswt_pff(weight_in_PopNB_mioi_oswt_pff)
    );
  SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp SysPE_PERun_weight_in_PopNB_mioi_weight_in_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .weight_in_PopNB_mioi_data_rsc_z_mxwt(weight_in_PopNB_mioi_data_rsc_z_mxwt),
      .weight_in_PopNB_mioi_return_rsc_z_mxwt(weight_in_PopNB_mioi_return_rsc_z_mxwt),
      .weight_in_PopNB_mioi_data_rsc_z(weight_in_PopNB_mioi_data_rsc_z),
      .weight_in_PopNB_mioi_biwt(weight_in_PopNB_mioi_biwt),
      .weight_in_PopNB_mioi_bdwt(weight_in_PopNB_mioi_bdwt),
      .weight_in_PopNB_mioi_return_rsc_z(weight_in_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_7_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_7_mioi (
  clk, rst, act_in_vec_7_val, act_in_vec_7_rdy, act_in_vec_7_msg, ReadRspRun_wen,
      act_in_vec_Push_7_mioi_oswt, act_in_vec_Push_7_mioi_wen_comp, act_in_vec_Push_7_mioi_m_rsc_dat_ReadRspRun,
      act_in_vec_Push_7_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_in_vec_7_val;
  input act_in_vec_7_rdy;
  output [7:0] act_in_vec_7_msg;
  input ReadRspRun_wen;
  input act_in_vec_Push_7_mioi_oswt;
  output act_in_vec_Push_7_mioi_wen_comp;
  input [7:0] act_in_vec_Push_7_mioi_m_rsc_dat_ReadRspRun;
  input act_in_vec_Push_7_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_in_vec_Push_7_mioi_biwt;
  wire act_in_vec_Push_7_mioi_bdwt;
  wire act_in_vec_Push_7_mioi_bcwt;
  wire act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  wire act_in_vec_Push_7_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_in_vec_Push_7_mioi
      (
      .this_val(act_in_vec_7_val),
      .this_rdy(act_in_vec_7_rdy),
      .this_msg(act_in_vec_7_msg),
      .m_rsc_dat(act_in_vec_Push_7_mioi_m_rsc_dat_ReadRspRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .ccs_ccore_done_sync_vld(act_in_vec_Push_7_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_act_in_vec_Push_7_mio_wait_ctrl InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_act_in_vec_Push_7_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_7_mioi_oswt(act_in_vec_Push_7_mioi_oswt),
      .act_in_vec_Push_7_mioi_biwt(act_in_vec_Push_7_mioi_biwt),
      .act_in_vec_Push_7_mioi_bdwt(act_in_vec_Push_7_mioi_bdwt),
      .act_in_vec_Push_7_mioi_bcwt(act_in_vec_Push_7_mioi_bcwt),
      .act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .act_in_vec_Push_7_mioi_ccs_ccore_done_sync_vld(act_in_vec_Push_7_mioi_ccs_ccore_done_sync_vld),
      .act_in_vec_Push_7_mioi_oswt_pff(act_in_vec_Push_7_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_act_in_vec_Push_7_mio_wait_dp InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_act_in_vec_Push_7_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_Push_7_mioi_oswt(act_in_vec_Push_7_mioi_oswt),
      .act_in_vec_Push_7_mioi_wen_comp(act_in_vec_Push_7_mioi_wen_comp),
      .act_in_vec_Push_7_mioi_biwt(act_in_vec_Push_7_mioi_biwt),
      .act_in_vec_Push_7_mioi_bdwt(act_in_vec_Push_7_mioi_bdwt),
      .act_in_vec_Push_7_mioi_bcwt(act_in_vec_Push_7_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_6_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_6_mioi (
  clk, rst, act_in_vec_6_val, act_in_vec_6_rdy, act_in_vec_6_msg, ReadRspRun_wen,
      act_in_vec_Push_6_mioi_oswt, act_in_vec_Push_6_mioi_wen_comp, act_in_vec_Push_6_mioi_m_rsc_dat_ReadRspRun,
      act_in_vec_Push_6_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_in_vec_6_val;
  input act_in_vec_6_rdy;
  output [7:0] act_in_vec_6_msg;
  input ReadRspRun_wen;
  input act_in_vec_Push_6_mioi_oswt;
  output act_in_vec_Push_6_mioi_wen_comp;
  input [7:0] act_in_vec_Push_6_mioi_m_rsc_dat_ReadRspRun;
  input act_in_vec_Push_6_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_in_vec_Push_6_mioi_biwt;
  wire act_in_vec_Push_6_mioi_bdwt;
  wire act_in_vec_Push_6_mioi_bcwt;
  wire act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  wire act_in_vec_Push_6_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_in_vec_Push_6_mioi
      (
      .this_val(act_in_vec_6_val),
      .this_rdy(act_in_vec_6_rdy),
      .this_msg(act_in_vec_6_msg),
      .m_rsc_dat(act_in_vec_Push_6_mioi_m_rsc_dat_ReadRspRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .ccs_ccore_done_sync_vld(act_in_vec_Push_6_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_act_in_vec_Push_6_mio_wait_ctrl InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_act_in_vec_Push_6_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_6_mioi_oswt(act_in_vec_Push_6_mioi_oswt),
      .act_in_vec_Push_6_mioi_biwt(act_in_vec_Push_6_mioi_biwt),
      .act_in_vec_Push_6_mioi_bdwt(act_in_vec_Push_6_mioi_bdwt),
      .act_in_vec_Push_6_mioi_bcwt(act_in_vec_Push_6_mioi_bcwt),
      .act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .act_in_vec_Push_6_mioi_ccs_ccore_done_sync_vld(act_in_vec_Push_6_mioi_ccs_ccore_done_sync_vld),
      .act_in_vec_Push_6_mioi_oswt_pff(act_in_vec_Push_6_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_act_in_vec_Push_6_mio_wait_dp InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_act_in_vec_Push_6_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_Push_6_mioi_oswt(act_in_vec_Push_6_mioi_oswt),
      .act_in_vec_Push_6_mioi_wen_comp(act_in_vec_Push_6_mioi_wen_comp),
      .act_in_vec_Push_6_mioi_biwt(act_in_vec_Push_6_mioi_biwt),
      .act_in_vec_Push_6_mioi_bdwt(act_in_vec_Push_6_mioi_bdwt),
      .act_in_vec_Push_6_mioi_bcwt(act_in_vec_Push_6_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_5_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_5_mioi (
  clk, rst, act_in_vec_5_val, act_in_vec_5_rdy, act_in_vec_5_msg, ReadRspRun_wen,
      act_in_vec_Push_5_mioi_oswt, act_in_vec_Push_5_mioi_wen_comp, act_in_vec_Push_5_mioi_m_rsc_dat_ReadRspRun,
      act_in_vec_Push_5_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_in_vec_5_val;
  input act_in_vec_5_rdy;
  output [7:0] act_in_vec_5_msg;
  input ReadRspRun_wen;
  input act_in_vec_Push_5_mioi_oswt;
  output act_in_vec_Push_5_mioi_wen_comp;
  input [7:0] act_in_vec_Push_5_mioi_m_rsc_dat_ReadRspRun;
  input act_in_vec_Push_5_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_in_vec_Push_5_mioi_biwt;
  wire act_in_vec_Push_5_mioi_bdwt;
  wire act_in_vec_Push_5_mioi_bcwt;
  wire act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  wire act_in_vec_Push_5_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_in_vec_Push_5_mioi
      (
      .this_val(act_in_vec_5_val),
      .this_rdy(act_in_vec_5_rdy),
      .this_msg(act_in_vec_5_msg),
      .m_rsc_dat(act_in_vec_Push_5_mioi_m_rsc_dat_ReadRspRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .ccs_ccore_done_sync_vld(act_in_vec_Push_5_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_act_in_vec_Push_5_mio_wait_ctrl InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_act_in_vec_Push_5_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_5_mioi_oswt(act_in_vec_Push_5_mioi_oswt),
      .act_in_vec_Push_5_mioi_biwt(act_in_vec_Push_5_mioi_biwt),
      .act_in_vec_Push_5_mioi_bdwt(act_in_vec_Push_5_mioi_bdwt),
      .act_in_vec_Push_5_mioi_bcwt(act_in_vec_Push_5_mioi_bcwt),
      .act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .act_in_vec_Push_5_mioi_ccs_ccore_done_sync_vld(act_in_vec_Push_5_mioi_ccs_ccore_done_sync_vld),
      .act_in_vec_Push_5_mioi_oswt_pff(act_in_vec_Push_5_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_act_in_vec_Push_5_mio_wait_dp InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_act_in_vec_Push_5_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_Push_5_mioi_oswt(act_in_vec_Push_5_mioi_oswt),
      .act_in_vec_Push_5_mioi_wen_comp(act_in_vec_Push_5_mioi_wen_comp),
      .act_in_vec_Push_5_mioi_biwt(act_in_vec_Push_5_mioi_biwt),
      .act_in_vec_Push_5_mioi_bdwt(act_in_vec_Push_5_mioi_bdwt),
      .act_in_vec_Push_5_mioi_bcwt(act_in_vec_Push_5_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_4_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_4_mioi (
  clk, rst, act_in_vec_4_val, act_in_vec_4_rdy, act_in_vec_4_msg, ReadRspRun_wen,
      act_in_vec_Push_4_mioi_oswt, act_in_vec_Push_4_mioi_wen_comp, act_in_vec_Push_4_mioi_m_rsc_dat_ReadRspRun,
      act_in_vec_Push_4_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_in_vec_4_val;
  input act_in_vec_4_rdy;
  output [7:0] act_in_vec_4_msg;
  input ReadRspRun_wen;
  input act_in_vec_Push_4_mioi_oswt;
  output act_in_vec_Push_4_mioi_wen_comp;
  input [7:0] act_in_vec_Push_4_mioi_m_rsc_dat_ReadRspRun;
  input act_in_vec_Push_4_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_in_vec_Push_4_mioi_biwt;
  wire act_in_vec_Push_4_mioi_bdwt;
  wire act_in_vec_Push_4_mioi_bcwt;
  wire act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  wire act_in_vec_Push_4_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_in_vec_Push_4_mioi
      (
      .this_val(act_in_vec_4_val),
      .this_rdy(act_in_vec_4_rdy),
      .this_msg(act_in_vec_4_msg),
      .m_rsc_dat(act_in_vec_Push_4_mioi_m_rsc_dat_ReadRspRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .ccs_ccore_done_sync_vld(act_in_vec_Push_4_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_act_in_vec_Push_4_mio_wait_ctrl InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_act_in_vec_Push_4_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_4_mioi_oswt(act_in_vec_Push_4_mioi_oswt),
      .act_in_vec_Push_4_mioi_biwt(act_in_vec_Push_4_mioi_biwt),
      .act_in_vec_Push_4_mioi_bdwt(act_in_vec_Push_4_mioi_bdwt),
      .act_in_vec_Push_4_mioi_bcwt(act_in_vec_Push_4_mioi_bcwt),
      .act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .act_in_vec_Push_4_mioi_ccs_ccore_done_sync_vld(act_in_vec_Push_4_mioi_ccs_ccore_done_sync_vld),
      .act_in_vec_Push_4_mioi_oswt_pff(act_in_vec_Push_4_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_act_in_vec_Push_4_mio_wait_dp InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_act_in_vec_Push_4_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_Push_4_mioi_oswt(act_in_vec_Push_4_mioi_oswt),
      .act_in_vec_Push_4_mioi_wen_comp(act_in_vec_Push_4_mioi_wen_comp),
      .act_in_vec_Push_4_mioi_biwt(act_in_vec_Push_4_mioi_biwt),
      .act_in_vec_Push_4_mioi_bdwt(act_in_vec_Push_4_mioi_bdwt),
      .act_in_vec_Push_4_mioi_bcwt(act_in_vec_Push_4_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_3_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_3_mioi (
  clk, rst, act_in_vec_3_val, act_in_vec_3_rdy, act_in_vec_3_msg, ReadRspRun_wen,
      act_in_vec_Push_3_mioi_oswt, act_in_vec_Push_3_mioi_wen_comp, act_in_vec_Push_3_mioi_m_rsc_dat_ReadRspRun,
      act_in_vec_Push_3_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_in_vec_3_val;
  input act_in_vec_3_rdy;
  output [7:0] act_in_vec_3_msg;
  input ReadRspRun_wen;
  input act_in_vec_Push_3_mioi_oswt;
  output act_in_vec_Push_3_mioi_wen_comp;
  input [7:0] act_in_vec_Push_3_mioi_m_rsc_dat_ReadRspRun;
  input act_in_vec_Push_3_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_in_vec_Push_3_mioi_biwt;
  wire act_in_vec_Push_3_mioi_bdwt;
  wire act_in_vec_Push_3_mioi_bcwt;
  wire act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  wire act_in_vec_Push_3_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_in_vec_Push_3_mioi
      (
      .this_val(act_in_vec_3_val),
      .this_rdy(act_in_vec_3_rdy),
      .this_msg(act_in_vec_3_msg),
      .m_rsc_dat(act_in_vec_Push_3_mioi_m_rsc_dat_ReadRspRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .ccs_ccore_done_sync_vld(act_in_vec_Push_3_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_act_in_vec_Push_3_mio_wait_ctrl InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_act_in_vec_Push_3_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_3_mioi_oswt(act_in_vec_Push_3_mioi_oswt),
      .act_in_vec_Push_3_mioi_biwt(act_in_vec_Push_3_mioi_biwt),
      .act_in_vec_Push_3_mioi_bdwt(act_in_vec_Push_3_mioi_bdwt),
      .act_in_vec_Push_3_mioi_bcwt(act_in_vec_Push_3_mioi_bcwt),
      .act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .act_in_vec_Push_3_mioi_ccs_ccore_done_sync_vld(act_in_vec_Push_3_mioi_ccs_ccore_done_sync_vld),
      .act_in_vec_Push_3_mioi_oswt_pff(act_in_vec_Push_3_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_act_in_vec_Push_3_mio_wait_dp InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_act_in_vec_Push_3_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_Push_3_mioi_oswt(act_in_vec_Push_3_mioi_oswt),
      .act_in_vec_Push_3_mioi_wen_comp(act_in_vec_Push_3_mioi_wen_comp),
      .act_in_vec_Push_3_mioi_biwt(act_in_vec_Push_3_mioi_biwt),
      .act_in_vec_Push_3_mioi_bdwt(act_in_vec_Push_3_mioi_bdwt),
      .act_in_vec_Push_3_mioi_bcwt(act_in_vec_Push_3_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_2_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_2_mioi (
  clk, rst, act_in_vec_2_val, act_in_vec_2_rdy, act_in_vec_2_msg, ReadRspRun_wen,
      act_in_vec_Push_2_mioi_oswt, act_in_vec_Push_2_mioi_wen_comp, act_in_vec_Push_2_mioi_m_rsc_dat_ReadRspRun,
      act_in_vec_Push_2_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_in_vec_2_val;
  input act_in_vec_2_rdy;
  output [7:0] act_in_vec_2_msg;
  input ReadRspRun_wen;
  input act_in_vec_Push_2_mioi_oswt;
  output act_in_vec_Push_2_mioi_wen_comp;
  input [7:0] act_in_vec_Push_2_mioi_m_rsc_dat_ReadRspRun;
  input act_in_vec_Push_2_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_in_vec_Push_2_mioi_biwt;
  wire act_in_vec_Push_2_mioi_bdwt;
  wire act_in_vec_Push_2_mioi_bcwt;
  wire act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  wire act_in_vec_Push_2_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_in_vec_Push_2_mioi
      (
      .this_val(act_in_vec_2_val),
      .this_rdy(act_in_vec_2_rdy),
      .this_msg(act_in_vec_2_msg),
      .m_rsc_dat(act_in_vec_Push_2_mioi_m_rsc_dat_ReadRspRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .ccs_ccore_done_sync_vld(act_in_vec_Push_2_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_act_in_vec_Push_2_mio_wait_ctrl InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_act_in_vec_Push_2_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_2_mioi_oswt(act_in_vec_Push_2_mioi_oswt),
      .act_in_vec_Push_2_mioi_biwt(act_in_vec_Push_2_mioi_biwt),
      .act_in_vec_Push_2_mioi_bdwt(act_in_vec_Push_2_mioi_bdwt),
      .act_in_vec_Push_2_mioi_bcwt(act_in_vec_Push_2_mioi_bcwt),
      .act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .act_in_vec_Push_2_mioi_ccs_ccore_done_sync_vld(act_in_vec_Push_2_mioi_ccs_ccore_done_sync_vld),
      .act_in_vec_Push_2_mioi_oswt_pff(act_in_vec_Push_2_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_act_in_vec_Push_2_mio_wait_dp InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_act_in_vec_Push_2_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_Push_2_mioi_oswt(act_in_vec_Push_2_mioi_oswt),
      .act_in_vec_Push_2_mioi_wen_comp(act_in_vec_Push_2_mioi_wen_comp),
      .act_in_vec_Push_2_mioi_biwt(act_in_vec_Push_2_mioi_biwt),
      .act_in_vec_Push_2_mioi_bdwt(act_in_vec_Push_2_mioi_bdwt),
      .act_in_vec_Push_2_mioi_bcwt(act_in_vec_Push_2_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_1_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_1_mioi (
  clk, rst, act_in_vec_1_val, act_in_vec_1_rdy, act_in_vec_1_msg, ReadRspRun_wen,
      act_in_vec_Push_1_mioi_oswt, act_in_vec_Push_1_mioi_wen_comp, act_in_vec_Push_1_mioi_m_rsc_dat_ReadRspRun,
      act_in_vec_Push_1_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_in_vec_1_val;
  input act_in_vec_1_rdy;
  output [7:0] act_in_vec_1_msg;
  input ReadRspRun_wen;
  input act_in_vec_Push_1_mioi_oswt;
  output act_in_vec_Push_1_mioi_wen_comp;
  input [7:0] act_in_vec_Push_1_mioi_m_rsc_dat_ReadRspRun;
  input act_in_vec_Push_1_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_in_vec_Push_1_mioi_biwt;
  wire act_in_vec_Push_1_mioi_bdwt;
  wire act_in_vec_Push_1_mioi_bcwt;
  wire act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  wire act_in_vec_Push_1_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_in_vec_Push_1_mioi
      (
      .this_val(act_in_vec_1_val),
      .this_rdy(act_in_vec_1_rdy),
      .this_msg(act_in_vec_1_msg),
      .m_rsc_dat(act_in_vec_Push_1_mioi_m_rsc_dat_ReadRspRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .ccs_ccore_done_sync_vld(act_in_vec_Push_1_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_act_in_vec_Push_1_mio_wait_ctrl InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_act_in_vec_Push_1_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_1_mioi_oswt(act_in_vec_Push_1_mioi_oswt),
      .act_in_vec_Push_1_mioi_biwt(act_in_vec_Push_1_mioi_biwt),
      .act_in_vec_Push_1_mioi_bdwt(act_in_vec_Push_1_mioi_bdwt),
      .act_in_vec_Push_1_mioi_bcwt(act_in_vec_Push_1_mioi_bcwt),
      .act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .act_in_vec_Push_1_mioi_ccs_ccore_done_sync_vld(act_in_vec_Push_1_mioi_ccs_ccore_done_sync_vld),
      .act_in_vec_Push_1_mioi_oswt_pff(act_in_vec_Push_1_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_act_in_vec_Push_1_mio_wait_dp InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_act_in_vec_Push_1_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_Push_1_mioi_oswt(act_in_vec_Push_1_mioi_oswt),
      .act_in_vec_Push_1_mioi_wen_comp(act_in_vec_Push_1_mioi_wen_comp),
      .act_in_vec_Push_1_mioi_biwt(act_in_vec_Push_1_mioi_biwt),
      .act_in_vec_Push_1_mioi_bdwt(act_in_vec_Push_1_mioi_bdwt),
      .act_in_vec_Push_1_mioi_bcwt(act_in_vec_Push_1_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_act_in_vec_Push_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_act_in_vec_Push_mioi (
  clk, rst, act_in_vec_0_val, act_in_vec_0_rdy, act_in_vec_0_msg, ReadRspRun_wen,
      act_in_vec_Push_mioi_oswt, act_in_vec_Push_mioi_wen_comp, act_in_vec_Push_mioi_m_rsc_dat_ReadRspRun,
      act_in_vec_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output act_in_vec_0_val;
  input act_in_vec_0_rdy;
  output [7:0] act_in_vec_0_msg;
  input ReadRspRun_wen;
  input act_in_vec_Push_mioi_oswt;
  output act_in_vec_Push_mioi_wen_comp;
  input [7:0] act_in_vec_Push_mioi_m_rsc_dat_ReadRspRun;
  input act_in_vec_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire act_in_vec_Push_mioi_biwt;
  wire act_in_vec_Push_mioi_bdwt;
  wire act_in_vec_Push_mioi_bcwt;
  wire act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;
  wire act_in_vec_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_OutBlocking_SysPE_InputType_Connections_SYN_PORT_Push  act_in_vec_Push_mioi
      (
      .this_val(act_in_vec_0_val),
      .this_rdy(act_in_vec_0_rdy),
      .this_msg(act_in_vec_0_msg),
      .m_rsc_dat(act_in_vec_Push_mioi_m_rsc_dat_ReadRspRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .ccs_ccore_done_sync_vld(act_in_vec_Push_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_mioi_act_in_vec_Push_mio_wait_ctrl InputSetup_ReadRspRun_act_in_vec_Push_mioi_act_in_vec_Push_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_mioi_oswt(act_in_vec_Push_mioi_oswt),
      .act_in_vec_Push_mioi_biwt(act_in_vec_Push_mioi_biwt),
      .act_in_vec_Push_mioi_bdwt(act_in_vec_Push_mioi_bdwt),
      .act_in_vec_Push_mioi_bcwt(act_in_vec_Push_mioi_bcwt),
      .act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .act_in_vec_Push_mioi_ccs_ccore_done_sync_vld(act_in_vec_Push_mioi_ccs_ccore_done_sync_vld),
      .act_in_vec_Push_mioi_oswt_pff(act_in_vec_Push_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_mioi_act_in_vec_Push_mio_wait_dp InputSetup_ReadRspRun_act_in_vec_Push_mioi_act_in_vec_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_Push_mioi_oswt(act_in_vec_Push_mioi_oswt),
      .act_in_vec_Push_mioi_wen_comp(act_in_vec_Push_mioi_wen_comp),
      .act_in_vec_Push_mioi_biwt(act_in_vec_Push_mioi_biwt),
      .act_in_vec_Push_mioi_bdwt(act_in_vec_Push_mioi_bdwt),
      .act_in_vec_Push_mioi_bcwt(act_in_vec_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun_rsp_inter_PopNB_mioi
// ------------------------------------------------------------------


module InputSetup_ReadRspRun_rsp_inter_PopNB_mioi (
  clk, rst, rsp_inter_val, rsp_inter_rdy, rsp_inter_msg, ReadRspRun_wen, rsp_inter_PopNB_mioi_oswt,
      ReadRspRun_wten, rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt, rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt,
      rsp_inter_PopNB_mioi_return_rsc_z_mxwt, rsp_inter_PopNB_mioi_oswt_pff
);
  input clk;
  input rst;
  input rsp_inter_val;
  output rsp_inter_rdy;
  input [71:0] rsp_inter_msg;
  input ReadRspRun_wen;
  input rsp_inter_PopNB_mioi_oswt;
  input ReadRspRun_wten;
  output [7:0] rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
  output [63:0] rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt;
  output rsp_inter_PopNB_mioi_return_rsc_z_mxwt;
  input rsp_inter_PopNB_mioi_oswt_pff;


  // Interconnect Declarations
  wire [7:0] rsp_inter_PopNB_mioi_data_valids_rsc_z;
  wire rsp_inter_PopNB_mioi_biwt;
  wire rsp_inter_PopNB_mioi_bdwt;
  wire [63:0] rsp_inter_PopNB_mioi_data_data_rsc_z;
  wire rsp_inter_PopNB_mioi_return_rsc_z;
  wire rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_PopNB
      rsp_inter_PopNB_mioi (
      .this_val(rsp_inter_val),
      .this_rdy(rsp_inter_rdy),
      .this_msg(rsp_inter_msg),
      .data_valids_rsc_z(rsp_inter_PopNB_mioi_data_valids_rsc_z),
      .data_data_rsc_z(rsp_inter_PopNB_mioi_data_data_rsc_z),
      .return_rsc_z(rsp_inter_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct)
    );
  InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_rsp_inter_PopNB_mio_wait_ctrl InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_rsp_inter_PopNB_mio_wait_ctrl_inst
      (
      .ReadRspRun_wen(ReadRspRun_wen),
      .rsp_inter_PopNB_mioi_oswt(rsp_inter_PopNB_mioi_oswt),
      .ReadRspRun_wten(ReadRspRun_wten),
      .rsp_inter_PopNB_mioi_biwt(rsp_inter_PopNB_mioi_biwt),
      .rsp_inter_PopNB_mioi_bdwt(rsp_inter_PopNB_mioi_bdwt),
      .rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct(rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_sct),
      .rsp_inter_PopNB_mioi_oswt_pff(rsp_inter_PopNB_mioi_oswt_pff)
    );
  InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_rsp_inter_PopNB_mio_wait_dp InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_rsp_inter_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt(rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt),
      .rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt(rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt),
      .rsp_inter_PopNB_mioi_return_rsc_z_mxwt(rsp_inter_PopNB_mioi_return_rsc_z_mxwt),
      .rsp_inter_PopNB_mioi_data_valids_rsc_z(rsp_inter_PopNB_mioi_data_valids_rsc_z),
      .rsp_inter_PopNB_mioi_biwt(rsp_inter_PopNB_mioi_biwt),
      .rsp_inter_PopNB_mioi_bdwt(rsp_inter_PopNB_mioi_bdwt),
      .rsp_inter_PopNB_mioi_data_data_rsc_z(rsp_inter_PopNB_mioi_data_data_rsc_z),
      .rsp_inter_PopNB_mioi_return_rsc_z(rsp_inter_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadReqRun_req_inter_PushNB_mioi
// ------------------------------------------------------------------


module InputSetup_ReadReqRun_req_inter_PushNB_mioi (
  clk, rst, req_inter_val, req_inter_rdy, req_inter_msg, req_inter_PushNB_mioi_m_valids_rsc_dat_ReadReqRun,
      req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff, req_inter_PushNB_mioi_iswt0_pff,
      ReadReqRun_wten_pff
);
  input clk;
  input rst;
  output req_inter_val;
  input req_inter_rdy;
  output [136:0] req_inter_msg;
  input [7:0] req_inter_PushNB_mioi_m_valids_rsc_dat_ReadReqRun;
  input [63:0] req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff;
  input req_inter_PushNB_mioi_iswt0_pff;
  input ReadReqRun_wten_pff;


  // Interconnect Declarations
  wire req_inter_PushNB_mioi_return_rsc_z;
  wire req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff;


  // Interconnect Declarations for Component Instantiations 
  wire [63:0] nl_req_inter_PushNB_mioi_m_addr_rsc_dat;
  assign nl_req_inter_PushNB_mioi_m_addr_rsc_dat = {(req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[63:49])
      , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff) , (req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[47:42])
      , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff) , (req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[40:34])
      , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff) , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff)
      , (req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[31:27]) , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff)
      , (req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[25:19]) , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff)
      , (req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[17]) , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff)
      , (req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[15:11]) , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff)
      , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff) , (req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[8:3])
      , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff) , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff)
      , (~ req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff)};
  Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PushNB
      req_inter_PushNB_mioi (
      .this_val(req_inter_val),
      .this_rdy(req_inter_rdy),
      .this_msg(req_inter_msg),
      .m_valids_rsc_dat(req_inter_PushNB_mioi_m_valids_rsc_dat_ReadReqRun),
      .m_addr_rsc_dat(nl_req_inter_PushNB_mioi_m_addr_rsc_dat[63:0]),
      .return_rsc_z(req_inter_PushNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff)
    );
  InputSetup_ReadReqRun_req_inter_PushNB_mioi_req_inter_PushNB_mio_wait_ctrl InputSetup_ReadReqRun_req_inter_PushNB_mioi_req_inter_PushNB_mio_wait_ctrl_inst
      (
      .req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_pff(req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_sct_iff),
      .req_inter_PushNB_mioi_iswt0_pff(req_inter_PushNB_mioi_iswt0_pff),
      .ReadReqRun_wten_pff(ReadReqRun_wten_pff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadReqRun_start_Pop_mioi
// ------------------------------------------------------------------


module InputSetup_ReadReqRun_start_Pop_mioi (
  clk, rst, start_val, start_rdy, start_msg, ReadReqRun_wen, start_Pop_mioi_return_rsc_z,
      start_Pop_mioi_oswt, ReadReqRun_wten, start_Pop_mioi_wen_comp, start_Pop_mioi_oswt_pff
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input [5:0] start_msg;
  input ReadReqRun_wen;
  output [5:0] start_Pop_mioi_return_rsc_z;
  input start_Pop_mioi_oswt;
  input ReadReqRun_wten;
  output start_Pop_mioi_wen_comp;
  input start_Pop_mioi_oswt_pff;


  // Interconnect Declarations
  wire start_Pop_mioi_biwt;
  wire start_Pop_mioi_bdwt;
  wire start_Pop_mioi_bcwt;
  wire start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_sct;
  wire start_Pop_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_InputSetup_StartType_Connections_SYN_PORT_Pop  start_Pop_mioi
      (
      .this_val(start_val),
      .this_rdy(start_rdy),
      .this_msg(start_msg),
      .return_rsc_z(start_Pop_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_sct),
      .ccs_ccore_done_sync_vld(start_Pop_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_ReadReqRun_start_Pop_mioi_start_Pop_mio_wait_ctrl InputSetup_ReadReqRun_start_Pop_mioi_start_Pop_mio_wait_ctrl_inst
      (
      .ReadReqRun_wen(ReadReqRun_wen),
      .start_Pop_mioi_oswt(start_Pop_mioi_oswt),
      .ReadReqRun_wten(ReadReqRun_wten),
      .start_Pop_mioi_biwt(start_Pop_mioi_biwt),
      .start_Pop_mioi_bdwt(start_Pop_mioi_bdwt),
      .start_Pop_mioi_bcwt(start_Pop_mioi_bcwt),
      .start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_sct(start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_sct),
      .start_Pop_mioi_ccs_ccore_done_sync_vld(start_Pop_mioi_ccs_ccore_done_sync_vld),
      .start_Pop_mioi_oswt_pff(start_Pop_mioi_oswt_pff)
    );
  InputSetup_ReadReqRun_start_Pop_mioi_start_Pop_mio_wait_dp InputSetup_ReadReqRun_start_Pop_mioi_start_Pop_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .start_Pop_mioi_oswt(start_Pop_mioi_oswt),
      .start_Pop_mioi_wen_comp(start_Pop_mioi_wen_comp),
      .start_Pop_mioi_biwt(start_Pop_mioi_biwt),
      .start_Pop_mioi_bdwt(start_Pop_mioi_bdwt),
      .start_Pop_mioi_bcwt(start_Pop_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_rsp_inter_Push_mioi
// ------------------------------------------------------------------


module InputSetup_MemoryRun_rsp_inter_Push_mioi (
  clk, rst, rsp_inter_val, rsp_inter_rdy, rsp_inter_msg, MemoryRun_wen, MemoryRun_wten,
      rsp_inter_Push_mioi_oswt, rsp_inter_Push_mioi_wen_comp, rsp_inter_Push_mioi_m_valids_rsc_dat_MemoryRun,
      rsp_inter_Push_mioi_m_data_rsc_dat_MemoryRun, rsp_inter_Push_mioi_oswt_pff
);
  input clk;
  input rst;
  output rsp_inter_val;
  input rsp_inter_rdy;
  output [71:0] rsp_inter_msg;
  input MemoryRun_wen;
  input MemoryRun_wten;
  input rsp_inter_Push_mioi_oswt;
  output rsp_inter_Push_mioi_wen_comp;
  input [7:0] rsp_inter_Push_mioi_m_valids_rsc_dat_MemoryRun;
  input [63:0] rsp_inter_Push_mioi_m_data_rsc_dat_MemoryRun;
  input rsp_inter_Push_mioi_oswt_pff;


  // Interconnect Declarations
  wire rsp_inter_Push_mioi_biwt;
  wire rsp_inter_Push_mioi_bdwt;
  wire rsp_inter_Push_mioi_bcwt;
  wire rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct;
  wire rsp_inter_Push_mioi_ccs_ccore_done_sync_vld;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_rsp_t_Connections_SYN_PORT_Push
      rsp_inter_Push_mioi (
      .this_val(rsp_inter_val),
      .this_rdy(rsp_inter_rdy),
      .this_msg(rsp_inter_msg),
      .m_valids_rsc_dat(rsp_inter_Push_mioi_m_valids_rsc_dat_MemoryRun),
      .m_data_rsc_dat(rsp_inter_Push_mioi_m_data_rsc_dat_MemoryRun),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct),
      .ccs_ccore_done_sync_vld(rsp_inter_Push_mioi_ccs_ccore_done_sync_vld)
    );
  InputSetup_MemoryRun_rsp_inter_Push_mioi_rsp_inter_Push_mio_wait_ctrl InputSetup_MemoryRun_rsp_inter_Push_mioi_rsp_inter_Push_mio_wait_ctrl_inst
      (
      .MemoryRun_wen(MemoryRun_wen),
      .MemoryRun_wten(MemoryRun_wten),
      .rsp_inter_Push_mioi_oswt(rsp_inter_Push_mioi_oswt),
      .rsp_inter_Push_mioi_biwt(rsp_inter_Push_mioi_biwt),
      .rsp_inter_Push_mioi_bdwt(rsp_inter_Push_mioi_bdwt),
      .rsp_inter_Push_mioi_bcwt(rsp_inter_Push_mioi_bcwt),
      .rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct(rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct),
      .rsp_inter_Push_mioi_ccs_ccore_done_sync_vld(rsp_inter_Push_mioi_ccs_ccore_done_sync_vld),
      .rsp_inter_Push_mioi_oswt_pff(rsp_inter_Push_mioi_oswt_pff)
    );
  InputSetup_MemoryRun_rsp_inter_Push_mioi_rsp_inter_Push_mio_wait_dp InputSetup_MemoryRun_rsp_inter_Push_mioi_rsp_inter_Push_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .rsp_inter_Push_mioi_oswt(rsp_inter_Push_mioi_oswt),
      .rsp_inter_Push_mioi_wen_comp(rsp_inter_Push_mioi_wen_comp),
      .rsp_inter_Push_mioi_biwt(rsp_inter_Push_mioi_biwt),
      .rsp_inter_Push_mioi_bdwt(rsp_inter_Push_mioi_bdwt),
      .rsp_inter_Push_mioi_bcwt(rsp_inter_Push_mioi_bcwt)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_write_req_PopNB_mioi
// ------------------------------------------------------------------


module InputSetup_MemoryRun_write_req_PopNB_mioi (
  clk, rst, write_req_val, write_req_rdy, write_req_msg, MemoryRun_wen, MemoryRun_wten,
      write_req_PopNB_mioi_oswt, write_req_PopNB_mioi_data_data_data_rsc_z_mxwt,
      write_req_PopNB_mioi_data_index_rsc_z_mxwt, write_req_PopNB_mioi_return_rsc_z_mxwt,
      write_req_PopNB_mioi_oswt_pff, MemoryRun_wten_pff
);
  input clk;
  input rst;
  input write_req_val;
  output write_req_rdy;
  input [68:0] write_req_msg;
  input MemoryRun_wen;
  input MemoryRun_wten;
  input write_req_PopNB_mioi_oswt;
  output [63:0] write_req_PopNB_mioi_data_data_data_rsc_z_mxwt;
  output [4:0] write_req_PopNB_mioi_data_index_rsc_z_mxwt;
  output write_req_PopNB_mioi_return_rsc_z_mxwt;
  input write_req_PopNB_mioi_oswt_pff;
  input MemoryRun_wten_pff;


  // Interconnect Declarations
  wire [63:0] write_req_PopNB_mioi_data_data_data_rsc_z;
  wire write_req_PopNB_mioi_biwt;
  wire write_req_PopNB_mioi_bdwt;
  wire [4:0] write_req_PopNB_mioi_data_index_rsc_z;
  wire write_req_PopNB_mioi_return_rsc_z;
  wire write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_InBlocking_InputSetup_WriteReq_Connections_SYN_PORT_PopNB  write_req_PopNB_mioi
      (
      .this_val(write_req_val),
      .this_rdy(write_req_rdy),
      .this_msg(write_req_msg),
      .data_data_data_rsc_z(write_req_PopNB_mioi_data_data_data_rsc_z),
      .data_index_rsc_z(write_req_PopNB_mioi_data_index_rsc_z),
      .return_rsc_z(write_req_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct)
    );
  InputSetup_MemoryRun_write_req_PopNB_mioi_write_req_PopNB_mio_wait_ctrl InputSetup_MemoryRun_write_req_PopNB_mioi_write_req_PopNB_mio_wait_ctrl_inst
      (
      .MemoryRun_wen(MemoryRun_wen),
      .MemoryRun_wten(MemoryRun_wten),
      .write_req_PopNB_mioi_oswt(write_req_PopNB_mioi_oswt),
      .write_req_PopNB_mioi_biwt(write_req_PopNB_mioi_biwt),
      .write_req_PopNB_mioi_bdwt(write_req_PopNB_mioi_bdwt),
      .write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct(write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct),
      .write_req_PopNB_mioi_oswt_pff(write_req_PopNB_mioi_oswt_pff),
      .MemoryRun_wten_pff(MemoryRun_wten_pff)
    );
  InputSetup_MemoryRun_write_req_PopNB_mioi_write_req_PopNB_mio_wait_dp InputSetup_MemoryRun_write_req_PopNB_mioi_write_req_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .write_req_PopNB_mioi_data_data_data_rsc_z_mxwt(write_req_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .write_req_PopNB_mioi_data_index_rsc_z_mxwt(write_req_PopNB_mioi_data_index_rsc_z_mxwt),
      .write_req_PopNB_mioi_return_rsc_z_mxwt(write_req_PopNB_mioi_return_rsc_z_mxwt),
      .write_req_PopNB_mioi_data_data_data_rsc_z(write_req_PopNB_mioi_data_data_data_rsc_z),
      .write_req_PopNB_mioi_biwt(write_req_PopNB_mioi_biwt),
      .write_req_PopNB_mioi_bdwt(write_req_PopNB_mioi_bdwt),
      .write_req_PopNB_mioi_data_index_rsc_z(write_req_PopNB_mioi_data_index_rsc_z),
      .write_req_PopNB_mioi_return_rsc_z(write_req_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun_req_inter_PopNB_mioi
// ------------------------------------------------------------------


module InputSetup_MemoryRun_req_inter_PopNB_mioi (
  clk, rst, req_inter_val, req_inter_rdy, req_inter_msg, MemoryRun_wen, req_inter_PopNB_mioi_oswt,
      MemoryRun_wten, req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt, req_inter_PopNB_mioi_data_valids_rsc_z_mxwt,
      req_inter_PopNB_mioi_data_addr_rsc_z_mxwt, req_inter_PopNB_mioi_data_data_rsc_z_mxwt,
      req_inter_PopNB_mioi_return_rsc_z_mxwt, req_inter_PopNB_mioi_oswt_pff, MemoryRun_wten_pff
);
  input clk;
  input rst;
  input req_inter_val;
  output req_inter_rdy;
  input [136:0] req_inter_msg;
  input MemoryRun_wen;
  input req_inter_PopNB_mioi_oswt;
  input MemoryRun_wten;
  output req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt;
  output [7:0] req_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
  output [63:0] req_inter_PopNB_mioi_data_addr_rsc_z_mxwt;
  output [63:0] req_inter_PopNB_mioi_data_data_rsc_z_mxwt;
  output req_inter_PopNB_mioi_return_rsc_z_mxwt;
  input req_inter_PopNB_mioi_oswt_pff;
  input MemoryRun_wten_pff;


  // Interconnect Declarations
  wire req_inter_PopNB_mioi_data_type_val_rsc_z;
  wire req_inter_PopNB_mioi_biwt;
  wire req_inter_PopNB_mioi_bdwt;
  wire [7:0] req_inter_PopNB_mioi_data_valids_rsc_z;
  wire [63:0] req_inter_PopNB_mioi_data_addr_rsc_z;
  wire [63:0] req_inter_PopNB_mioi_data_data_rsc_z;
  wire req_inter_PopNB_mioi_return_rsc_z;
  wire req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_ArbitratedScratchpad_InputSetup_InputType_256U_8U_8U_0U_req_t_Connections_SYN_PORT_PopNB
      req_inter_PopNB_mioi (
      .this_val(req_inter_val),
      .this_rdy(req_inter_rdy),
      .this_msg(req_inter_msg),
      .data_type_val_rsc_z(req_inter_PopNB_mioi_data_type_val_rsc_z),
      .data_valids_rsc_z(req_inter_PopNB_mioi_data_valids_rsc_z),
      .data_addr_rsc_z(req_inter_PopNB_mioi_data_addr_rsc_z),
      .data_data_rsc_z(req_inter_PopNB_mioi_data_data_rsc_z),
      .return_rsc_z(req_inter_PopNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct)
    );
  InputSetup_MemoryRun_req_inter_PopNB_mioi_req_inter_PopNB_mio_wait_ctrl InputSetup_MemoryRun_req_inter_PopNB_mioi_req_inter_PopNB_mio_wait_ctrl_inst
      (
      .MemoryRun_wen(MemoryRun_wen),
      .req_inter_PopNB_mioi_oswt(req_inter_PopNB_mioi_oswt),
      .MemoryRun_wten(MemoryRun_wten),
      .req_inter_PopNB_mioi_biwt(req_inter_PopNB_mioi_biwt),
      .req_inter_PopNB_mioi_bdwt(req_inter_PopNB_mioi_bdwt),
      .req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct(req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_sct),
      .req_inter_PopNB_mioi_oswt_pff(req_inter_PopNB_mioi_oswt_pff),
      .MemoryRun_wten_pff(MemoryRun_wten_pff)
    );
  InputSetup_MemoryRun_req_inter_PopNB_mioi_req_inter_PopNB_mio_wait_dp InputSetup_MemoryRun_req_inter_PopNB_mioi_req_inter_PopNB_mio_wait_dp_inst
      (
      .clk(clk),
      .rst(rst),
      .req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt(req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt),
      .req_inter_PopNB_mioi_data_valids_rsc_z_mxwt(req_inter_PopNB_mioi_data_valids_rsc_z_mxwt),
      .req_inter_PopNB_mioi_data_addr_rsc_z_mxwt(req_inter_PopNB_mioi_data_addr_rsc_z_mxwt),
      .req_inter_PopNB_mioi_data_data_rsc_z_mxwt(req_inter_PopNB_mioi_data_data_rsc_z_mxwt),
      .req_inter_PopNB_mioi_return_rsc_z_mxwt(req_inter_PopNB_mioi_return_rsc_z_mxwt),
      .req_inter_PopNB_mioi_data_type_val_rsc_z(req_inter_PopNB_mioi_data_type_val_rsc_z),
      .req_inter_PopNB_mioi_biwt(req_inter_PopNB_mioi_biwt),
      .req_inter_PopNB_mioi_bdwt(req_inter_PopNB_mioi_bdwt),
      .req_inter_PopNB_mioi_data_valids_rsc_z(req_inter_PopNB_mioi_data_valids_rsc_z),
      .req_inter_PopNB_mioi_data_addr_rsc_z(req_inter_PopNB_mioi_data_addr_rsc_z),
      .req_inter_PopNB_mioi_data_data_rsc_z(req_inter_PopNB_mioi_data_data_rsc_z),
      .req_inter_PopNB_mioi_return_rsc_z(req_inter_PopNB_mioi_return_rsc_z)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE_PERun
// ------------------------------------------------------------------


module SysPE_PERun (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, act_in_val, act_in_rdy,
      act_in_msg, accum_in_val, accum_in_rdy, accum_in_msg, act_out_val, act_out_rdy,
      act_out_msg, accum_out_val, accum_out_rdy, accum_out_msg, weight_out_val, weight_out_rdy,
      weight_out_msg
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;


  // Interconnect Declarations
  wire PERun_wen;
  wire PERun_wten;
  wire [7:0] weight_in_PopNB_mioi_data_rsc_z_mxwt;
  wire weight_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [7:0] act_in_PopNB_mioi_data_rsc_z_mxwt;
  wire act_in_PopNB_mioi_return_rsc_z_mxwt;
  wire [31:0] accum_in_PopNB_mioi_data_rsc_z_mxwt;
  wire accum_in_PopNB_mioi_return_rsc_z_mxwt;
  wire act_out_Push_mioi_wen_comp;
  wire accum_out_Push_mioi_wen_comp;
  wire [1:0] fsm_output;
  wire while_while_or_tmp;
  wire is_accum_in_sva_dfm_1;
  reg is_accum_in_sva;
  reg while_stage_0_3;
  reg is_act_in_sva;
  wire while_land_lpi_1_dfm_1;
  reg reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  reg reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  wire is_accum_in_63_and_cse;
  wire and_1_cse;
  wire and_8_rmff;
  wire and_7_rmff;
  reg [7:0] weight_reg_sva;
  reg [7:0] act_reg_sva;
  wire [7:0] act_out_Push_mioi_m_rsc_dat_PERun_mx1;
  wire [31:0] accum_reg_sva_mx0;
  reg [31:0] accum_reg_sva;

  wire[0:0] mux_7_nl;
  wire[0:0] or_10_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] or_12_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] nor_1_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] nor_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff;
  assign nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff =
      fsm_output[1];
  wire [0:0] nl_SysPE_PERun_weight_out_PushNB_mioi_inst_PERun_wten;
  assign nl_SysPE_PERun_weight_out_PushNB_mioi_inst_PERun_wten = ~ PERun_wen;
  wire [0:0] nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_iswt0;
  assign nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_iswt0
      = weight_in_PopNB_mioi_return_rsc_z_mxwt & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  wire [7:0] nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_m_rsc_dat_PERun;
  assign nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_m_rsc_dat_PERun
      = weight_reg_sva;
  wire[0:0] act_reg_63_and_1_nl;
  wire [7:0] nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun;
  assign act_reg_63_and_1_nl = (~ is_act_in_sva) & (fsm_output[1]);
  assign nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun
      = MUX_v_8_2_2(act_reg_sva, act_in_PopNB_mioi_data_rsc_z_mxwt, act_reg_63_and_1_nl);
  wire[15:0] while_if_3_accum_out_reg_mul_nl;
  wire [31:0] nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun;
  assign while_if_3_accum_out_reg_mul_nl = conv_s2u_16_16($signed((act_out_Push_mioi_m_rsc_dat_PERun_mx1))
      * $signed(weight_reg_sva));
  assign nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun
      = conv_s2u_16_32(while_if_3_accum_out_reg_mul_nl) + accum_reg_sva_mx0;
  SysPE_PERun_weight_in_PopNB_mioi SysPE_PERun_weight_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_val),
      .weight_in_rdy(weight_in_rdy),
      .weight_in_msg(weight_in_msg),
      .PERun_wen(PERun_wen),
      .weight_in_PopNB_mioi_oswt(reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .PERun_wten(PERun_wten),
      .weight_in_PopNB_mioi_data_rsc_z_mxwt(weight_in_PopNB_mioi_data_rsc_z_mxwt),
      .weight_in_PopNB_mioi_return_rsc_z_mxwt(weight_in_PopNB_mioi_return_rsc_z_mxwt),
      .weight_in_PopNB_mioi_oswt_pff(nl_SysPE_PERun_weight_in_PopNB_mioi_inst_weight_in_PopNB_mioi_oswt_pff[0:0])
    );
  SysPE_PERun_weight_out_PushNB_mioi SysPE_PERun_weight_out_PushNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .weight_out_val(weight_out_val),
      .weight_out_rdy(weight_out_rdy),
      .weight_out_msg(weight_out_msg),
      .PERun_wten(nl_SysPE_PERun_weight_out_PushNB_mioi_inst_PERun_wten[0:0]),
      .weight_out_PushNB_mioi_iswt0(nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_iswt0[0:0]),
      .weight_out_PushNB_mioi_m_rsc_dat_PERun(nl_SysPE_PERun_weight_out_PushNB_mioi_inst_weight_out_PushNB_mioi_m_rsc_dat_PERun[7:0])
    );
  SysPE_PERun_act_in_PopNB_mioi SysPE_PERun_act_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .act_in_val(act_in_val),
      .act_in_rdy(act_in_rdy),
      .act_in_msg(act_in_msg),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_in_PopNB_mioi_oswt(reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .act_in_PopNB_mioi_data_rsc_z_mxwt(act_in_PopNB_mioi_data_rsc_z_mxwt),
      .act_in_PopNB_mioi_return_rsc_z_mxwt(act_in_PopNB_mioi_return_rsc_z_mxwt),
      .act_in_PopNB_mioi_oswt_pff(and_8_rmff)
    );
  SysPE_PERun_accum_in_PopNB_mioi SysPE_PERun_accum_in_PopNB_mioi_inst (
      .clk(clk),
      .rst(rst),
      .accum_in_val(accum_in_val),
      .accum_in_rdy(accum_in_rdy),
      .accum_in_msg(accum_in_msg),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .accum_in_PopNB_mioi_oswt(reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .accum_in_PopNB_mioi_data_rsc_z_mxwt(accum_in_PopNB_mioi_data_rsc_z_mxwt),
      .accum_in_PopNB_mioi_return_rsc_z_mxwt(accum_in_PopNB_mioi_return_rsc_z_mxwt),
      .accum_in_PopNB_mioi_oswt_pff(and_7_rmff)
    );
  SysPE_PERun_act_out_Push_mioi SysPE_PERun_act_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .act_out_val(act_out_val),
      .act_out_rdy(act_out_rdy),
      .act_out_msg(act_out_msg),
      .PERun_wen(PERun_wen),
      .act_out_Push_mioi_oswt(reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .act_out_Push_mioi_m_rsc_dat_PERun(nl_SysPE_PERun_act_out_Push_mioi_inst_act_out_Push_mioi_m_rsc_dat_PERun[7:0]),
      .act_out_Push_mioi_oswt_pff(and_1_cse)
    );
  SysPE_PERun_accum_out_Push_mioi SysPE_PERun_accum_out_Push_mioi_inst (
      .clk(clk),
      .rst(rst),
      .accum_out_val(accum_out_val),
      .accum_out_rdy(accum_out_rdy),
      .accum_out_msg(accum_out_msg),
      .PERun_wen(PERun_wen),
      .accum_out_Push_mioi_oswt(reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_m_rsc_dat_PERun(nl_SysPE_PERun_accum_out_Push_mioi_inst_accum_out_Push_mioi_m_rsc_dat_PERun[31:0]),
      .accum_out_Push_mioi_oswt_pff(and_1_cse)
    );
  SysPE_PERun_staller SysPE_PERun_staller_inst (
      .clk(clk),
      .rst(rst),
      .PERun_wen(PERun_wen),
      .PERun_wten(PERun_wten),
      .act_out_Push_mioi_wen_comp(act_out_Push_mioi_wen_comp),
      .accum_out_Push_mioi_wen_comp(accum_out_Push_mioi_wen_comp)
    );
  SysPE_PERun_PERun_fsm SysPE_PERun_PERun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .PERun_wen(PERun_wen),
      .fsm_output(fsm_output)
    );
  assign and_1_cse = while_while_or_tmp & is_accum_in_sva_dfm_1 & while_stage_0_3;
  assign or_10_nl = (~ is_accum_in_sva_dfm_1) | act_in_PopNB_mioi_return_rsc_z_mxwt
      | is_act_in_sva;
  assign mux_7_nl = MUX_s_1_2_2((~ is_accum_in_sva), (or_10_nl), while_stage_0_3);
  assign and_7_rmff = (mux_7_nl) & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  assign or_12_nl = is_accum_in_sva_dfm_1 | (~ while_while_or_tmp);
  assign mux_8_nl = MUX_s_1_2_2((~ is_act_in_sva), (or_12_nl), while_stage_0_3);
  assign and_8_rmff = (mux_8_nl) & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
  assign is_accum_in_63_and_cse = PERun_wen & while_stage_0_3;
  assign act_out_Push_mioi_m_rsc_dat_PERun_mx1 = MUX_v_8_2_2(act_in_PopNB_mioi_data_rsc_z_mxwt,
      act_reg_sva, is_act_in_sva);
  assign accum_reg_sva_mx0 = MUX_v_32_2_2(accum_in_PopNB_mioi_data_rsc_z_mxwt, accum_reg_sva,
      is_accum_in_sva);
  assign is_accum_in_sva_dfm_1 = accum_in_PopNB_mioi_return_rsc_z_mxwt | is_accum_in_sva;
  assign while_land_lpi_1_dfm_1 = is_accum_in_sva_dfm_1 & while_while_or_tmp;
  assign while_while_or_tmp = act_in_PopNB_mioi_return_rsc_z_mxwt | is_act_in_sva;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= 1'b0;
      while_stage_0_3 <= 1'b0;
    end
    else if ( PERun_wen ) begin
      reg_accum_out_Push_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_1_cse;
      reg_accum_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_7_rmff;
      reg_act_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= and_8_rmff;
      reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse <= fsm_output[1];
      while_stage_0_3 <= reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      is_accum_in_sva <= 1'b0;
      is_act_in_sva <= 1'b0;
    end
    else if ( is_accum_in_63_and_cse ) begin
      is_accum_in_sva <= is_accum_in_sva_dfm_1 & (~ while_land_lpi_1_dfm_1);
      is_act_in_sva <= while_while_or_tmp & (~ while_land_lpi_1_dfm_1);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      weight_reg_sva <= 8'b00000000;
    end
    else if ( PERun_wen & weight_in_PopNB_mioi_return_rsc_z_mxwt & reg_weight_in_PopNB_mioi_ccs_ccore_start_rsc_dat_PERun_psct_cse
        ) begin
      weight_reg_sva <= weight_in_PopNB_mioi_data_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      accum_reg_sva <= 32'b00000000000000000000000000000000;
    end
    else if ( PERun_wen & (mux_5_nl) ) begin
      accum_reg_sva <= accum_reg_sva_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      act_reg_sva <= 8'b00000000;
    end
    else if ( PERun_wen & (mux_6_nl) ) begin
      act_reg_sva <= act_out_Push_mioi_m_rsc_dat_PERun_mx1;
    end
  end
  assign nor_1_nl = ~((~ is_accum_in_sva_dfm_1) | act_in_PopNB_mioi_return_rsc_z_mxwt
      | is_act_in_sva);
  assign mux_5_nl = MUX_s_1_2_2(is_accum_in_sva, (nor_1_nl), while_stage_0_3);
  assign nor_nl = ~(is_accum_in_sva_dfm_1 | (~ while_while_or_tmp));
  assign mux_6_nl = MUX_s_1_2_2(is_act_in_sva, (nor_nl), while_stage_0_3);

  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [31:0] MUX_v_32_2_2;
    input [31:0] input_0;
    input [31:0] input_1;
    input [0:0] sel;
    reg [31:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_32_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [15:0] conv_s2u_16_16 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_16 = vector;
  end
  endfunction


  function automatic [31:0] conv_s2u_16_32 ;
    input [15:0]  vector ;
  begin
    conv_s2u_16_32 = {{16{vector[15]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadRspRun
// ------------------------------------------------------------------


module InputSetup_ReadRspRun (
  clk, rst, act_in_vec_0_val, act_in_vec_1_val, act_in_vec_2_val, act_in_vec_3_val,
      act_in_vec_4_val, act_in_vec_5_val, act_in_vec_6_val, act_in_vec_7_val, act_in_vec_0_rdy,
      act_in_vec_1_rdy, act_in_vec_2_rdy, act_in_vec_3_rdy, act_in_vec_4_rdy, act_in_vec_5_rdy,
      act_in_vec_6_rdy, act_in_vec_7_rdy, act_in_vec_0_msg, act_in_vec_1_msg, act_in_vec_2_msg,
      act_in_vec_3_msg, act_in_vec_4_msg, act_in_vec_5_msg, act_in_vec_6_msg, act_in_vec_7_msg,
      rsp_inter_val, rsp_inter_rdy, rsp_inter_msg
);
  input clk;
  input rst;
  output act_in_vec_0_val;
  output act_in_vec_1_val;
  output act_in_vec_2_val;
  output act_in_vec_3_val;
  output act_in_vec_4_val;
  output act_in_vec_5_val;
  output act_in_vec_6_val;
  output act_in_vec_7_val;
  input act_in_vec_0_rdy;
  input act_in_vec_1_rdy;
  input act_in_vec_2_rdy;
  input act_in_vec_3_rdy;
  input act_in_vec_4_rdy;
  input act_in_vec_5_rdy;
  input act_in_vec_6_rdy;
  input act_in_vec_7_rdy;
  output [7:0] act_in_vec_0_msg;
  output [7:0] act_in_vec_1_msg;
  output [7:0] act_in_vec_2_msg;
  output [7:0] act_in_vec_3_msg;
  output [7:0] act_in_vec_4_msg;
  output [7:0] act_in_vec_5_msg;
  output [7:0] act_in_vec_6_msg;
  output [7:0] act_in_vec_7_msg;
  input rsp_inter_val;
  output rsp_inter_rdy;
  input [71:0] rsp_inter_msg;


  // Interconnect Declarations
  wire ReadRspRun_wen;
  wire ReadRspRun_wten;
  wire [7:0] rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
  wire [63:0] rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt;
  wire rsp_inter_PopNB_mioi_return_rsc_z_mxwt;
  wire act_in_vec_Push_mioi_wen_comp;
  wire act_in_vec_Push_1_mioi_wen_comp;
  wire act_in_vec_Push_2_mioi_wen_comp;
  wire act_in_vec_Push_3_mioi_wen_comp;
  wire act_in_vec_Push_4_mioi_wen_comp;
  wire act_in_vec_Push_5_mioi_wen_comp;
  wire act_in_vec_Push_6_mioi_wen_comp;
  wire act_in_vec_Push_7_mioi_wen_comp;
  wire [1:0] fsm_output;
  wire and_dcpl;
  reg reg_act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  reg reg_act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  reg reg_act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  reg reg_act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  reg reg_act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  reg reg_act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  reg reg_act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  reg reg_act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  reg reg_rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  wire and_8_rmff;
  wire and_7_rmff;
  wire and_6_rmff;
  wire and_5_rmff;
  wire and_4_rmff;
  wire and_3_rmff;
  wire and_2_rmff;
  wire and_1_rmff;

  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_1;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_2;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_3;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_4;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_5;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_6;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_prb_7;
  wire[0:0] p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_inst_rsp_inter_PopNB_mioi_oswt_pff;
  assign nl_InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_inst_rsp_inter_PopNB_mioi_oswt_pff
      = fsm_output[1];
  wire [7:0] nl_InputSetup_ReadRspRun_act_in_vec_Push_mioi_inst_act_in_vec_Push_mioi_m_rsc_dat_ReadRspRun;
  assign nl_InputSetup_ReadRspRun_act_in_vec_Push_mioi_inst_act_in_vec_Push_mioi_m_rsc_dat_ReadRspRun
      = rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt[7:0];
  wire [7:0] nl_InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_inst_act_in_vec_Push_1_mioi_m_rsc_dat_ReadRspRun;
  assign nl_InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_inst_act_in_vec_Push_1_mioi_m_rsc_dat_ReadRspRun
      = rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt[15:8];
  wire [7:0] nl_InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_inst_act_in_vec_Push_2_mioi_m_rsc_dat_ReadRspRun;
  assign nl_InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_inst_act_in_vec_Push_2_mioi_m_rsc_dat_ReadRspRun
      = rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt[23:16];
  wire [7:0] nl_InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_inst_act_in_vec_Push_3_mioi_m_rsc_dat_ReadRspRun;
  assign nl_InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_inst_act_in_vec_Push_3_mioi_m_rsc_dat_ReadRspRun
      = rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt[31:24];
  wire [7:0] nl_InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_inst_act_in_vec_Push_4_mioi_m_rsc_dat_ReadRspRun;
  assign nl_InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_inst_act_in_vec_Push_4_mioi_m_rsc_dat_ReadRspRun
      = rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt[39:32];
  wire [7:0] nl_InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_inst_act_in_vec_Push_5_mioi_m_rsc_dat_ReadRspRun;
  assign nl_InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_inst_act_in_vec_Push_5_mioi_m_rsc_dat_ReadRspRun
      = rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt[47:40];
  wire [7:0] nl_InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_inst_act_in_vec_Push_6_mioi_m_rsc_dat_ReadRspRun;
  assign nl_InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_inst_act_in_vec_Push_6_mioi_m_rsc_dat_ReadRspRun
      = rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt[55:48];
  wire [7:0] nl_InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_inst_act_in_vec_Push_7_mioi_m_rsc_dat_ReadRspRun;
  assign nl_InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_inst_act_in_vec_Push_7_mioi_m_rsc_dat_ReadRspRun
      = rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt[63:56];
  InputSetup_ReadRspRun_rsp_inter_PopNB_mioi InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rsp_inter_val(rsp_inter_val),
      .rsp_inter_rdy(rsp_inter_rdy),
      .rsp_inter_msg(rsp_inter_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .rsp_inter_PopNB_mioi_oswt(reg_rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .ReadRspRun_wten(ReadRspRun_wten),
      .rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt(rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt),
      .rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt(rsp_inter_PopNB_mioi_data_data_rsc_z_mxwt),
      .rsp_inter_PopNB_mioi_return_rsc_z_mxwt(rsp_inter_PopNB_mioi_return_rsc_z_mxwt),
      .rsp_inter_PopNB_mioi_oswt_pff(nl_InputSetup_ReadRspRun_rsp_inter_PopNB_mioi_inst_rsp_inter_PopNB_mioi_oswt_pff[0:0])
    );
  InputSetup_ReadRspRun_act_in_vec_Push_mioi InputSetup_ReadRspRun_act_in_vec_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_0_val(act_in_vec_0_val),
      .act_in_vec_0_rdy(act_in_vec_0_rdy),
      .act_in_vec_0_msg(act_in_vec_0_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_mioi_oswt(reg_act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .act_in_vec_Push_mioi_wen_comp(act_in_vec_Push_mioi_wen_comp),
      .act_in_vec_Push_mioi_m_rsc_dat_ReadRspRun(nl_InputSetup_ReadRspRun_act_in_vec_Push_mioi_inst_act_in_vec_Push_mioi_m_rsc_dat_ReadRspRun[7:0]),
      .act_in_vec_Push_mioi_oswt_pff(and_8_rmff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_1_mioi InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_1_val(act_in_vec_1_val),
      .act_in_vec_1_rdy(act_in_vec_1_rdy),
      .act_in_vec_1_msg(act_in_vec_1_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_1_mioi_oswt(reg_act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .act_in_vec_Push_1_mioi_wen_comp(act_in_vec_Push_1_mioi_wen_comp),
      .act_in_vec_Push_1_mioi_m_rsc_dat_ReadRspRun(nl_InputSetup_ReadRspRun_act_in_vec_Push_1_mioi_inst_act_in_vec_Push_1_mioi_m_rsc_dat_ReadRspRun[7:0]),
      .act_in_vec_Push_1_mioi_oswt_pff(and_7_rmff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_2_mioi InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_2_val(act_in_vec_2_val),
      .act_in_vec_2_rdy(act_in_vec_2_rdy),
      .act_in_vec_2_msg(act_in_vec_2_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_2_mioi_oswt(reg_act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .act_in_vec_Push_2_mioi_wen_comp(act_in_vec_Push_2_mioi_wen_comp),
      .act_in_vec_Push_2_mioi_m_rsc_dat_ReadRspRun(nl_InputSetup_ReadRspRun_act_in_vec_Push_2_mioi_inst_act_in_vec_Push_2_mioi_m_rsc_dat_ReadRspRun[7:0]),
      .act_in_vec_Push_2_mioi_oswt_pff(and_6_rmff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_3_mioi InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_3_val(act_in_vec_3_val),
      .act_in_vec_3_rdy(act_in_vec_3_rdy),
      .act_in_vec_3_msg(act_in_vec_3_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_3_mioi_oswt(reg_act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .act_in_vec_Push_3_mioi_wen_comp(act_in_vec_Push_3_mioi_wen_comp),
      .act_in_vec_Push_3_mioi_m_rsc_dat_ReadRspRun(nl_InputSetup_ReadRspRun_act_in_vec_Push_3_mioi_inst_act_in_vec_Push_3_mioi_m_rsc_dat_ReadRspRun[7:0]),
      .act_in_vec_Push_3_mioi_oswt_pff(and_5_rmff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_4_mioi InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_4_val(act_in_vec_4_val),
      .act_in_vec_4_rdy(act_in_vec_4_rdy),
      .act_in_vec_4_msg(act_in_vec_4_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_4_mioi_oswt(reg_act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .act_in_vec_Push_4_mioi_wen_comp(act_in_vec_Push_4_mioi_wen_comp),
      .act_in_vec_Push_4_mioi_m_rsc_dat_ReadRspRun(nl_InputSetup_ReadRspRun_act_in_vec_Push_4_mioi_inst_act_in_vec_Push_4_mioi_m_rsc_dat_ReadRspRun[7:0]),
      .act_in_vec_Push_4_mioi_oswt_pff(and_4_rmff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_5_mioi InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_5_val(act_in_vec_5_val),
      .act_in_vec_5_rdy(act_in_vec_5_rdy),
      .act_in_vec_5_msg(act_in_vec_5_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_5_mioi_oswt(reg_act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .act_in_vec_Push_5_mioi_wen_comp(act_in_vec_Push_5_mioi_wen_comp),
      .act_in_vec_Push_5_mioi_m_rsc_dat_ReadRspRun(nl_InputSetup_ReadRspRun_act_in_vec_Push_5_mioi_inst_act_in_vec_Push_5_mioi_m_rsc_dat_ReadRspRun[7:0]),
      .act_in_vec_Push_5_mioi_oswt_pff(and_3_rmff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_6_mioi InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_6_val(act_in_vec_6_val),
      .act_in_vec_6_rdy(act_in_vec_6_rdy),
      .act_in_vec_6_msg(act_in_vec_6_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_6_mioi_oswt(reg_act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .act_in_vec_Push_6_mioi_wen_comp(act_in_vec_Push_6_mioi_wen_comp),
      .act_in_vec_Push_6_mioi_m_rsc_dat_ReadRspRun(nl_InputSetup_ReadRspRun_act_in_vec_Push_6_mioi_inst_act_in_vec_Push_6_mioi_m_rsc_dat_ReadRspRun[7:0]),
      .act_in_vec_Push_6_mioi_oswt_pff(and_2_rmff)
    );
  InputSetup_ReadRspRun_act_in_vec_Push_7_mioi InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .act_in_vec_7_val(act_in_vec_7_val),
      .act_in_vec_7_rdy(act_in_vec_7_rdy),
      .act_in_vec_7_msg(act_in_vec_7_msg),
      .ReadRspRun_wen(ReadRspRun_wen),
      .act_in_vec_Push_7_mioi_oswt(reg_act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse),
      .act_in_vec_Push_7_mioi_wen_comp(act_in_vec_Push_7_mioi_wen_comp),
      .act_in_vec_Push_7_mioi_m_rsc_dat_ReadRspRun(nl_InputSetup_ReadRspRun_act_in_vec_Push_7_mioi_inst_act_in_vec_Push_7_mioi_m_rsc_dat_ReadRspRun[7:0]),
      .act_in_vec_Push_7_mioi_oswt_pff(and_1_rmff)
    );
  InputSetup_ReadRspRun_staller_2 InputSetup_ReadRspRun_staller_2_inst (
      .clk(clk),
      .rst(rst),
      .ReadRspRun_wen(ReadRspRun_wen),
      .ReadRspRun_wten(ReadRspRun_wten),
      .act_in_vec_Push_mioi_wen_comp(act_in_vec_Push_mioi_wen_comp),
      .act_in_vec_Push_1_mioi_wen_comp(act_in_vec_Push_1_mioi_wen_comp),
      .act_in_vec_Push_2_mioi_wen_comp(act_in_vec_Push_2_mioi_wen_comp),
      .act_in_vec_Push_3_mioi_wen_comp(act_in_vec_Push_3_mioi_wen_comp),
      .act_in_vec_Push_4_mioi_wen_comp(act_in_vec_Push_4_mioi_wen_comp),
      .act_in_vec_Push_5_mioi_wen_comp(act_in_vec_Push_5_mioi_wen_comp),
      .act_in_vec_Push_6_mioi_wen_comp(act_in_vec_Push_6_mioi_wen_comp),
      .act_in_vec_Push_7_mioi_wen_comp(act_in_vec_Push_7_mioi_wen_comp)
    );
  InputSetup_ReadRspRun_ReadRspRun_fsm InputSetup_ReadRspRun_ReadRspRun_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .ReadRspRun_wen(ReadRspRun_wen),
      .fsm_output(fsm_output)
    );
  assign p0_Unreachable_virtual_function_in_abstract_class_prb = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 2309
  // psl default clock = (posedge clk);
  // psl InputSetup_ReadRspRun_connections_h_ln2309_assert_0_and_Unreachablevirtualfunctioninabstractclassnot : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb  -> p0_Unreachable_virtual_function_in_abstract_class_prb );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_1 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 2309
  // psl default clock = (posedge clk);
  // psl InputSetup_ReadRspRun_connections_h_ln2309_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_1 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1  -> p0_Unreachable_virtual_function_in_abstract_class_prb_1 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_1 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_2 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 2309
  // psl default clock = (posedge clk);
  // psl InputSetup_ReadRspRun_connections_h_ln2309_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_2 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2  -> p0_Unreachable_virtual_function_in_abstract_class_prb_2 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_2 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_3 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 2309
  // psl default clock = (posedge clk);
  // psl InputSetup_ReadRspRun_connections_h_ln2309_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_3 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3  -> p0_Unreachable_virtual_function_in_abstract_class_prb_3 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_3 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_4 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 2309
  // psl default clock = (posedge clk);
  // psl InputSetup_ReadRspRun_connections_h_ln2309_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_4 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4  -> p0_Unreachable_virtual_function_in_abstract_class_prb_4 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_4 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_5 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 2309
  // psl default clock = (posedge clk);
  // psl InputSetup_ReadRspRun_connections_h_ln2309_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_5 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5  -> p0_Unreachable_virtual_function_in_abstract_class_prb_5 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_5 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_6 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 2309
  // psl default clock = (posedge clk);
  // psl InputSetup_ReadRspRun_connections_h_ln2309_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_6 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6  -> p0_Unreachable_virtual_function_in_abstract_class_prb_6 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_6 = 1'b0;
  assign p0_Unreachable_virtual_function_in_abstract_class_prb_7 = 1'b0;
  // assert(0 && "Unreachable virtual function in abstract class!") - ../../../matchlib/connections/include/connections/connections.h: line 2309
  // psl default clock = (posedge clk);
  // psl InputSetup_ReadRspRun_connections_h_ln2309_assert_0_and_Unreachablevirtualfunctioninabstractclassnot_7 : assert always ( rst &&  p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7  -> p0_Unreachable_virtual_function_in_abstract_class_prb_7 );
  assign p0_Unreachable_virtual_function_in_abstract_class_ctrl_prb_7 = 1'b0;
  assign and_1_rmff = and_dcpl & (rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt[7]);
  assign and_2_rmff = and_dcpl & (rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt[6]);
  assign and_3_rmff = and_dcpl & (rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt[5]);
  assign and_4_rmff = and_dcpl & (rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt[4]);
  assign and_5_rmff = and_dcpl & (rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt[3]);
  assign and_6_rmff = and_dcpl & (rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt[2]);
  assign and_7_rmff = and_dcpl & (rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt[1]);
  assign and_8_rmff = and_dcpl & (rsp_inter_PopNB_mioi_data_valids_rsc_z_mxwt[0]);
  assign and_dcpl = rsp_inter_PopNB_mioi_return_rsc_z_mxwt & reg_rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse;
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
      reg_act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
      reg_act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
      reg_act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
      reg_act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
      reg_act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
      reg_act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
      reg_act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
      reg_rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= 1'b0;
    end
    else if ( ReadRspRun_wen ) begin
      reg_act_in_vec_Push_7_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= and_1_rmff;
      reg_act_in_vec_Push_6_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= and_2_rmff;
      reg_act_in_vec_Push_5_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= and_3_rmff;
      reg_act_in_vec_Push_4_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= and_4_rmff;
      reg_act_in_vec_Push_3_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= and_5_rmff;
      reg_act_in_vec_Push_2_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= and_6_rmff;
      reg_act_in_vec_Push_1_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= and_7_rmff;
      reg_act_in_vec_Push_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= and_8_rmff;
      reg_rsp_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_ReadRspRun_psct_cse <= fsm_output[1];
    end
  end
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_ReadReqRun
// ------------------------------------------------------------------


module InputSetup_ReadReqRun (
  clk, rst, start_val, start_rdy, start_msg, req_inter_val, req_inter_rdy, req_inter_msg
);
  input clk;
  input rst;
  input start_val;
  output start_rdy;
  input [5:0] start_msg;
  output req_inter_val;
  input req_inter_rdy;
  output [136:0] req_inter_msg;


  // Interconnect Declarations
  wire [5:0] start_Pop_mioi_return_rsc_z;
  wire start_Pop_mioi_wen_comp;
  wire [5:0] fsm_output;
  wire or_tmp_7;
  reg exit_while_if_for_sva;
  wire operator_6_false_slc_operator_6_false_acc_7_svs_mx1;
  wire [7:0] operator_6_false_acc_2_cse_1;
  wire [8:0] nl_operator_6_false_acc_2_cse_1;
  reg [5:0] while_M_sva;
  reg [6:0] while_if_for_t_7_0_sva_6_0;
  reg reg_start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_psct_cse;
  wire ReadReqRun_wten_iff;
  wire while_if_for_if_for_mux_1_rmff;
  wire while_if_for_if_for_mux_rmff;
  wire while_req_reg_addr_mux_2_rmff;
  wire while_if_for_t_mux_rmff;
  wire while_req_reg_addr_mux_rmff;
  wire while_if_for_if_for_mux_2_rmff;
  wire while_req_reg_addr_mux_1_rmff;
  wire [4:0] while_if_for_else_if_for_6_if_conc_1_pmx_7_3_lpi_2_dfm_1;
  wire while_if_for_asn_37;
  wire while_if_for_asn_39;
  wire [3:0] while_if_for_else_if_for_3_if_conc_1_pmx_7_4_lpi_2_dfm_1;
  wire while_if_for_else_while_if_for_else_or_9_cse;
  wire while_if_for_else_while_if_for_else_or_8_cse;
  wire while_if_for_else_while_if_for_else_or_10_cse;
  wire [3:0] z_out;
  wire [4:0] nl_z_out;
  wire [3:0] z_out_1;
  wire [4:0] nl_z_out_1;
  wire [4:0] z_out_2;
  wire [5:0] nl_z_out_2;
  wire [4:0] z_out_3;
  wire [5:0] nl_z_out_3;
  wire [4:0] z_out_4;
  wire [5:0] nl_z_out_4;
  wire [3:0] z_out_5;
  wire [4:0] nl_z_out_5;
  wire [4:0] z_out_6;
  wire [5:0] nl_z_out_6;
  wire [7:0] z_out_7;
  wire [8:0] nl_z_out_7;
  reg [6:0] operator_33_true_return_6_0_sva;
  reg operator_6_false_slc_operator_6_false_acc_7_svs;
  wire and_33_cse;
  wire and_37_cse;
  wire operator_6_false_acc_itm_7_1;
  wire operator_6_false_acc_12_itm_6;
  wire operator_6_false_acc_11_itm_7_1;
  wire operator_6_false_acc_9_itm_7_1;
  wire operator_6_false_acc_10_itm_5;
  wire operator_6_false_acc_8_itm_6_1;
  wire while_if_for_else_if_for_2_operator_6_false_acc_itm_7_1;
  wire while_if_for_if_acc_itm_4_1;
  wire [1:0] while_if_for_if_for_if_while_if_for_if_for_if_and_cse;
  wire [5:0] z_out_8_7_2;

  wire[0:0] while_if_for_else_while_if_for_else_or_7_nl;
  wire[0:0] while_if_for_else_while_if_for_else_or_3_nl;
  wire[0:0] while_if_for_else_while_if_for_else_or_4_nl;
  wire[0:0] while_if_for_else_while_if_for_else_or_6_nl;
  wire[8:0] while_if_for_acc_nl;
  wire[10:0] nl_while_if_for_acc_nl;
  wire[6:0] while_if_for_t_mux_1_nl;
  wire[0:0] not_nl;
  wire[7:0] operator_6_false_acc_nl;
  wire[9:0] nl_operator_6_false_acc_nl;
  wire[6:0] operator_6_false_acc_12_nl;
  wire[7:0] nl_operator_6_false_acc_12_nl;
  wire[7:0] operator_6_false_acc_11_nl;
  wire[8:0] nl_operator_6_false_acc_11_nl;
  wire[7:0] operator_6_false_acc_9_nl;
  wire[8:0] nl_operator_6_false_acc_9_nl;
  wire[5:0] operator_6_false_acc_10_nl;
  wire[6:0] nl_operator_6_false_acc_10_nl;
  wire[6:0] operator_6_false_acc_8_nl;
  wire[7:0] nl_operator_6_false_acc_8_nl;
  wire[7:0] while_if_for_else_if_for_2_operator_6_false_acc_nl;
  wire[8:0] nl_while_if_for_else_if_for_2_operator_6_false_acc_nl;
  wire[4:0] while_if_for_if_acc_nl;
  wire[5:0] nl_while_if_for_if_acc_nl;
  wire[2:0] while_if_for_if_for_if_mux_11_nl;
  wire[3:0] while_if_for_else_if_for_if_mux_5_nl;
  wire[1:0] while_if_for_if_for_if_while_if_for_if_for_if_or_1_nl;
  wire[0:0] not_42_nl;
  wire[1:0] while_if_for_else_if_for_if_mux_6_nl;
  wire[6:0] operator_6_false_mux_1_nl;
  wire[7:0] while_if_for_if_for_if_acc_nl;
  wire[8:0] nl_while_if_for_if_for_if_acc_nl;
  wire[7:0] while_if_for_if_for_if_mux_12_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_InputSetup_ReadReqRun_start_Pop_mioi_inst_start_Pop_mioi_oswt_pff;
  assign nl_InputSetup_ReadReqRun_start_Pop_mioi_inst_start_Pop_mioi_oswt_pff = fsm_output[1];
  wire[0:0] while_if_for_while_if_for_or_nl;
  wire [7:0] nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_m_valids_rsc_dat_ReadReqRun;
  assign while_if_for_while_if_for_or_nl = operator_6_false_acc_itm_7_1 | operator_6_false_slc_operator_6_false_acc_7_svs_mx1
      | while_if_for_if_acc_itm_4_1;
  assign nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_m_valids_rsc_dat_ReadReqRun
      = {while_if_for_if_for_mux_1_rmff , while_if_for_if_for_mux_rmff , while_req_reg_addr_mux_2_rmff
      , while_if_for_t_mux_rmff , while_req_reg_addr_mux_rmff , while_if_for_if_for_mux_2_rmff
      , while_req_reg_addr_mux_1_rmff , (while_if_for_while_if_for_or_nl)};
  wire[4:0] and_28_nl;
  wire[4:0] mux_2_nl;
  wire[0:0] and_nl;
  wire[0:0] nor_nl;
  wire[3:0] and_29_nl;
  wire[3:0] mux_3_nl;
  wire[0:0] and_19_nl;
  wire[0:0] nor_7_nl;
  wire[0:0] while_if_for_if_for_mux_4_nl;
  wire[0:0] while_if_for_else_mux_38_nl;
  wire[0:0] while_if_for_else_if_for_while_if_for_else_if_for_and_9_nl;
  wire[0:0] while_if_for_if_for_while_if_for_if_for_and_8_nl;
  wire[3:0] while_if_for_while_if_for_mux1h_5_nl;
  wire[0:0] while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_3_nl;
  wire[0:0] while_if_for_while_if_for_mux1h_3_nl;
  wire[0:0] while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_2_nl;
  wire[2:0] and_30_nl;
  wire[2:0] mux_4_nl;
  wire[0:0] and_21_nl;
  wire[0:0] nor_8_nl;
  wire[1:0] mux_9_nl;
  wire[1:0] and_31_nl;
  wire[0:0] nor_9_nl;
  wire[0:0] and_68_nl;
  wire[4:0] mux_nl;
  wire[3:0] while_if_for_while_if_for_while_if_for_mux_nl;
  wire[2:0] while_if_for_if_for_while_if_for_if_for_and_3_nl;
  wire[0:0] while_if_for_if_for_not_13_nl;
  wire[0:0] or_19_nl;
  wire[2:0] while_if_for_while_if_for_mux1h_6_nl;
  wire[0:0] while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_1_nl;
  wire[0:0] while_if_for_while_if_for_mux1h_1_nl;
  wire[0:0] while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_nl;
  wire[0:0] while_if_for_if_for_mux_3_nl;
  wire[0:0] while_if_for_else_mux_37_nl;
  wire[0:0] while_if_for_else_if_for_while_if_for_else_if_for_and_3_nl;
  wire[0:0] while_if_for_if_for_while_if_for_if_for_and_7_nl;
  wire[4:0] mux_1_nl;
  wire[3:0] while_if_for_while_if_for_while_if_for_mux_1_nl;
  wire[2:0] while_if_for_if_for_while_if_for_if_for_and_nl;
  wire[0:0] while_if_for_if_for_not_8_nl;
  wire[0:0] or_20_nl;
  wire[1:0] while_if_for_while_if_for_and_nl;
  wire[2:0] while_if_for_while_if_for_and_4_nl;
  wire[0:0] while_if_for_or_nl;
  wire [63:0] nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff;
  assign and_nl = while_if_for_else_while_if_for_else_or_9_cse & (~ while_if_for_if_acc_itm_4_1);
  assign mux_2_nl = MUX_v_5_2_2((signext_5_1(~ operator_6_false_acc_itm_7_1)), z_out_3,
      and_nl);
  assign nor_nl = ~((~(operator_6_false_acc_itm_7_1 | operator_6_false_acc_12_itm_6))
      | while_if_for_if_acc_itm_4_1);
  assign and_28_nl = MUX_v_5_2_2(5'b00000, (mux_2_nl), (nor_nl));
  assign and_19_nl = while_if_for_else_while_if_for_else_or_8_cse & (~ while_if_for_if_acc_itm_4_1);
  assign mux_3_nl = MUX_v_4_2_2((signext_4_1(~ operator_6_false_acc_itm_7_1)), z_out_1,
      and_19_nl);
  assign nor_7_nl = ~((~(operator_6_false_acc_itm_7_1 | operator_6_false_acc_11_itm_7_1))
      | while_if_for_if_acc_itm_4_1);
  assign and_29_nl = MUX_v_4_2_2(4'b0000, (mux_3_nl), (nor_7_nl));
  assign while_if_for_else_if_for_while_if_for_else_if_for_and_9_nl = (while_if_for_t_7_0_sva_6_0[0])
      & operator_6_false_acc_11_itm_7_1;
  assign while_if_for_else_mux_38_nl = MUX_s_1_2_2((while_if_for_else_if_for_while_if_for_else_if_for_and_9_nl),
      (while_if_for_t_7_0_sva_6_0[0]), operator_6_false_acc_itm_7_1);
  assign while_if_for_if_for_while_if_for_if_for_and_8_nl = (while_if_for_t_7_0_sva_6_0[0])
      & (~ (z_out_8_7_2[0]));
  assign while_if_for_if_for_mux_4_nl = MUX_s_1_2_2((while_if_for_else_mux_38_nl),
      (while_if_for_if_for_while_if_for_if_for_and_8_nl), while_if_for_if_acc_itm_4_1);
  assign while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_3_nl = ~(((while_if_for_t_7_0_sva_6_0[0])
      ^ (while_if_for_t_7_0_sva_6_0[1])) | (z_out[3]));
  assign while_if_for_while_if_for_mux1h_5_nl = MUX1HOT_v_4_3_2((while_if_for_else_if_for_6_if_conc_1_pmx_7_3_lpi_2_dfm_1[4:1]),
      (z_out_4[4:1]), ({3'b000 , (while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_3_nl)}),
      {while_if_for_asn_37 , while_if_for_asn_39 , while_if_for_if_acc_itm_4_1});
  assign while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_2_nl = ~((while_if_for_t_7_0_sva_6_0[0])
      | (z_out[3]));
  assign while_if_for_while_if_for_mux1h_3_nl = MUX1HOT_s_1_3_2((while_if_for_else_if_for_6_if_conc_1_pmx_7_3_lpi_2_dfm_1[0]),
      (z_out_4[0]), (while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_2_nl),
      {while_if_for_asn_37 , while_if_for_asn_39 , while_if_for_if_acc_itm_4_1});
  assign and_21_nl = while_if_for_else_while_if_for_else_or_10_cse & (~ while_if_for_if_acc_itm_4_1);
  assign mux_4_nl = MUX_v_3_2_2((signext_3_1(~ operator_6_false_acc_itm_7_1)), (z_out[2:0]),
      and_21_nl);
  assign nor_8_nl = ~((~(operator_6_false_acc_itm_7_1 | operator_6_false_acc_9_itm_7_1))
      | while_if_for_if_acc_itm_4_1);
  assign and_30_nl = MUX_v_3_2_2(3'b000, (mux_4_nl), (nor_8_nl));
  assign nor_9_nl = ~((while_if_for_if_acc_itm_4_1 & (~ (while_if_for_t_7_0_sva_6_0[2])))
      | (while_if_for_asn_37 & (~ operator_6_false_acc_9_itm_7_1)));
  assign and_31_nl = MUX_v_2_2_2(2'b00, (signext_2_1(nor_9_nl)), while_if_for_asn_37);
  assign and_68_nl = ((while_if_for_t_7_0_sva_6_0[2]) | (~ while_if_for_if_acc_itm_4_1))
      & (operator_6_false_acc_9_itm_7_1 | (~ while_if_for_asn_37));
  assign mux_9_nl = MUX_v_2_2_2((and_31_nl), (while_if_for_t_7_0_sva_6_0[1:0]), and_68_nl);
  assign while_if_for_if_for_not_13_nl = ~ (z_out_6[3]);
  assign while_if_for_if_for_while_if_for_if_for_and_3_nl = MUX_v_3_2_2(3'b000, (z_out_1[2:0]),
      (while_if_for_if_for_not_13_nl));
  assign while_if_for_while_if_for_while_if_for_mux_nl = MUX_v_4_2_2(({{3{operator_6_false_acc_8_itm_6_1}},
      operator_6_false_acc_8_itm_6_1}), ({1'b0 , (while_if_for_if_for_while_if_for_if_for_and_3_nl)}),
      while_if_for_if_acc_itm_4_1);
  assign or_19_nl = (while_if_for_asn_37 & operator_6_false_acc_8_itm_6_1) | while_if_for_asn_39;
  assign mux_nl = MUX_v_5_2_2((signext_5_4(while_if_for_while_if_for_while_if_for_mux_nl)),
      z_out_2, or_19_nl);
  assign while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_1_nl = ~(((while_if_for_t_7_0_sva_6_0[1])
      ^ (while_if_for_t_7_0_sva_6_0[2])) | (z_out_5[2]));
  assign while_if_for_while_if_for_mux1h_6_nl = MUX1HOT_v_3_3_2((while_if_for_else_if_for_3_if_conc_1_pmx_7_4_lpi_2_dfm_1[3:1]),
      (z_out_5[3:1]), ({2'b00 , (while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_1_nl)}),
      {while_if_for_asn_37 , while_if_for_asn_39 , while_if_for_if_acc_itm_4_1});
  assign while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_nl = ~((while_if_for_t_7_0_sva_6_0[1])
      | (z_out_5[2]));
  assign while_if_for_while_if_for_mux1h_1_nl = MUX1HOT_s_1_3_2((while_if_for_else_if_for_3_if_conc_1_pmx_7_4_lpi_2_dfm_1[0]),
      (z_out_5[0]), (while_if_for_if_for_while_if_for_if_for_while_if_for_if_for_nor_nl),
      {while_if_for_asn_37 , while_if_for_asn_39 , while_if_for_if_acc_itm_4_1});
  assign while_if_for_else_if_for_while_if_for_else_if_for_and_3_nl = (while_if_for_t_7_0_sva_6_0[0])
      & (z_out_8_7_2[5]);
  assign while_if_for_else_mux_37_nl = MUX_s_1_2_2((while_if_for_else_if_for_while_if_for_else_if_for_and_3_nl),
      (while_if_for_t_7_0_sva_6_0[0]), operator_6_false_acc_itm_7_1);
  assign while_if_for_if_for_while_if_for_if_for_and_7_nl = (while_if_for_t_7_0_sva_6_0[0])
      & (~ (z_out_5[2]));
  assign while_if_for_if_for_mux_3_nl = MUX_s_1_2_2((while_if_for_else_mux_37_nl),
      (while_if_for_if_for_while_if_for_if_for_and_7_nl), while_if_for_if_acc_itm_4_1);
  assign while_if_for_if_for_not_8_nl = ~ (z_out_3[3]);
  assign while_if_for_if_for_while_if_for_if_for_and_nl = MUX_v_3_2_2(3'b000, (z_out_4[2:0]),
      (while_if_for_if_for_not_8_nl));
  assign while_if_for_while_if_for_while_if_for_mux_1_nl = MUX_v_4_2_2(({{3{while_if_for_else_if_for_2_operator_6_false_acc_itm_7_1}},
      while_if_for_else_if_for_2_operator_6_false_acc_itm_7_1}), ({1'b0 , (while_if_for_if_for_while_if_for_if_for_and_nl)}),
      while_if_for_if_acc_itm_4_1);
  assign or_20_nl = (while_if_for_asn_37 & while_if_for_else_if_for_2_operator_6_false_acc_itm_7_1)
      | while_if_for_asn_39;
  assign mux_1_nl = MUX_v_5_2_2((signext_5_4(while_if_for_while_if_for_while_if_for_mux_1_nl)),
      z_out_6, or_20_nl);
  assign while_if_for_while_if_for_and_nl = (while_if_for_t_7_0_sva_6_0[4:3]) & ({{1{operator_6_false_slc_operator_6_false_acc_7_svs_mx1}},
      operator_6_false_slc_operator_6_false_acc_7_svs_mx1}) & (signext_2_1(~ while_if_for_if_acc_itm_4_1));
  assign while_if_for_or_nl = operator_6_false_slc_operator_6_false_acc_7_svs_mx1
      | while_if_for_if_acc_itm_4_1;
  assign while_if_for_while_if_for_and_4_nl = MUX_v_3_2_2(3'b000, (while_if_for_t_7_0_sva_6_0[2:0]),
      (while_if_for_or_nl));
  assign nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff
      = {(and_28_nl) , ({{2{while_if_for_if_for_mux_1_rmff}}, while_if_for_if_for_mux_1_rmff})
      , (and_29_nl) , (while_if_for_if_for_mux_4_nl) , ({{1{while_if_for_if_for_mux_rmff}},
      while_if_for_if_for_mux_rmff}) , 1'b0 , (while_if_for_while_if_for_mux1h_5_nl)
      , (while_if_for_while_if_for_mux1h_3_nl) , while_req_reg_addr_mux_2_rmff ,
      1'b0 , while_req_reg_addr_mux_2_rmff , (and_30_nl) , (mux_9_nl) , while_if_for_t_mux_rmff
      , 2'b00 , (mux_nl) , 1'b0 , ({{1{while_req_reg_addr_mux_rmff}}, while_req_reg_addr_mux_rmff})
      , (while_if_for_while_if_for_mux1h_6_nl) , (while_if_for_while_if_for_mux1h_1_nl)
      , (while_if_for_if_for_mux_3_nl) , 1'b0 , while_if_for_if_for_mux_2_rmff ,
      1'b0 , (mux_1_nl) , 2'b00 , while_req_reg_addr_mux_1_rmff , (while_if_for_while_if_for_and_nl)
      , (while_if_for_while_if_for_and_4_nl) , 3'b000};
  wire [0:0] nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_iswt0_pff;
  assign nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_iswt0_pff
      = fsm_output[3];
  wire [0:0] nl_InputSetup_ReadReqRun_ReadReqRun_fsm_inst_while_C_1_tr0;
  assign nl_InputSetup_ReadReqRun_ReadReqRun_fsm_inst_while_C_1_tr0 = ~((start_Pop_mioi_return_rsc_z!=6'b000000));
  InputSetup_ReadReqRun_start_Pop_mioi InputSetup_ReadReqRun_start_Pop_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .ReadReqRun_wen(start_Pop_mioi_wen_comp),
      .start_Pop_mioi_return_rsc_z(start_Pop_mioi_return_rsc_z),
      .start_Pop_mioi_oswt(reg_start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_psct_cse),
      .ReadReqRun_wten(ReadReqRun_wten_iff),
      .start_Pop_mioi_wen_comp(start_Pop_mioi_wen_comp),
      .start_Pop_mioi_oswt_pff(nl_InputSetup_ReadReqRun_start_Pop_mioi_inst_start_Pop_mioi_oswt_pff[0:0])
    );
  InputSetup_ReadReqRun_req_inter_PushNB_mioi InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .req_inter_val(req_inter_val),
      .req_inter_rdy(req_inter_rdy),
      .req_inter_msg(req_inter_msg),
      .req_inter_PushNB_mioi_m_valids_rsc_dat_ReadReqRun(nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_m_valids_rsc_dat_ReadReqRun[7:0]),
      .req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff(nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_m_addr_rsc_dat_ReadReqRun_pff[63:0]),
      .req_inter_PushNB_mioi_iswt0_pff(nl_InputSetup_ReadReqRun_req_inter_PushNB_mioi_inst_req_inter_PushNB_mioi_iswt0_pff[0:0]),
      .ReadReqRun_wten_pff(ReadReqRun_wten_iff)
    );
  InputSetup_ReadReqRun_staller_1 InputSetup_ReadReqRun_staller_1_inst (
      .start_Pop_mioi_wen_comp(start_Pop_mioi_wen_comp),
      .ReadReqRun_wten_pff(ReadReqRun_wten_iff)
    );
  InputSetup_ReadReqRun_ReadReqRun_fsm InputSetup_ReadReqRun_ReadReqRun_fsm_inst
      (
      .clk(clk),
      .rst(rst),
      .start_Pop_mioi_wen_comp(start_Pop_mioi_wen_comp),
      .fsm_output(fsm_output),
      .while_C_1_tr0(nl_InputSetup_ReadReqRun_ReadReqRun_fsm_inst_while_C_1_tr0[0:0]),
      .while_if_for_C_1_tr0(exit_while_if_for_sva)
    );
  assign while_if_for_else_while_if_for_else_or_7_nl = operator_6_false_acc_8_itm_6_1
      | operator_6_false_acc_itm_7_1;
  assign while_req_reg_addr_mux_rmff = MUX_s_1_2_2((while_if_for_else_while_if_for_else_or_7_nl),
      (~ (z_out_6[3])), while_if_for_if_acc_itm_4_1);
  assign while_if_for_else_while_if_for_else_or_8_cse = operator_6_false_acc_11_itm_7_1
      | operator_6_false_acc_itm_7_1;
  assign while_if_for_if_for_mux_rmff = MUX_s_1_2_2(while_if_for_else_while_if_for_else_or_8_cse,
      (~ (z_out_8_7_2[0])), while_if_for_if_acc_itm_4_1);
  assign while_if_for_else_while_if_for_else_or_9_cse = operator_6_false_acc_12_itm_6
      | operator_6_false_acc_itm_7_1;
  assign while_if_for_if_for_mux_1_rmff = MUX_s_1_2_2(while_if_for_else_while_if_for_else_or_9_cse,
      (~ (z_out_2[3])), while_if_for_if_acc_itm_4_1);
  assign while_if_for_else_while_if_for_else_or_3_nl = while_if_for_else_if_for_2_operator_6_false_acc_itm_7_1
      | operator_6_false_acc_itm_7_1;
  assign while_req_reg_addr_mux_1_rmff = MUX_s_1_2_2((while_if_for_else_while_if_for_else_or_3_nl),
      (~ (z_out_3[3])), while_if_for_if_acc_itm_4_1);
  assign while_if_for_else_while_if_for_else_or_4_nl = (z_out_8_7_2[5]) | operator_6_false_acc_itm_7_1;
  assign while_if_for_if_for_mux_2_rmff = MUX_s_1_2_2((while_if_for_else_while_if_for_else_or_4_nl),
      (~ (z_out_5[2])), while_if_for_if_acc_itm_4_1);
  assign while_if_for_else_while_if_for_else_or_10_cse = operator_6_false_acc_9_itm_7_1
      | operator_6_false_acc_itm_7_1;
  assign while_if_for_t_mux_rmff = MUX_s_1_2_2(while_if_for_else_while_if_for_else_or_10_cse,
      (while_if_for_t_7_0_sva_6_0[2]), while_if_for_if_acc_itm_4_1);
  assign while_if_for_else_while_if_for_else_or_6_nl = operator_6_false_acc_10_itm_5
      | operator_6_false_acc_itm_7_1;
  assign while_req_reg_addr_mux_2_rmff = MUX_s_1_2_2((while_if_for_else_while_if_for_else_or_6_nl),
      (~ (z_out[3])), while_if_for_if_acc_itm_4_1);
  assign nl_operator_6_false_acc_nl = conv_u2s_7_8(while_if_for_t_7_0_sva_6_0) +
      conv_s2s_7_8({1'b1 , (~ while_M_sva)}) + 8'b00000001;
  assign operator_6_false_acc_nl = nl_operator_6_false_acc_nl[7:0];
  assign operator_6_false_acc_itm_7_1 = readslicef_8_1_7((operator_6_false_acc_nl));
  assign operator_6_false_slc_operator_6_false_acc_7_svs_mx1 = MUX_s_1_2_2(operator_6_false_acc_itm_7_1,
      operator_6_false_slc_operator_6_false_acc_7_svs, while_if_for_if_acc_itm_4_1);
  assign nl_operator_6_false_acc_12_nl = (operator_6_false_acc_2_cse_1[7:1]) + 7'b1011101;
  assign operator_6_false_acc_12_nl = nl_operator_6_false_acc_12_nl[6:0];
  assign operator_6_false_acc_12_itm_6 = readslicef_7_1_6((operator_6_false_acc_12_nl));
  assign nl_operator_6_false_acc_11_nl = operator_6_false_acc_2_cse_1 + 8'b10111011;
  assign operator_6_false_acc_11_nl = nl_operator_6_false_acc_11_nl[7:0];
  assign operator_6_false_acc_11_itm_7_1 = readslicef_8_1_7((operator_6_false_acc_11_nl));
  assign while_if_for_else_if_for_6_if_conc_1_pmx_7_3_lpi_2_dfm_1 = MUX_v_5_2_2(5'b00000,
      z_out_4, operator_6_false_acc_10_itm_5);
  assign nl_operator_6_false_acc_9_nl = operator_6_false_acc_2_cse_1 + 8'b10111101;
  assign operator_6_false_acc_9_nl = nl_operator_6_false_acc_9_nl[7:0];
  assign operator_6_false_acc_9_itm_7_1 = readslicef_8_1_7((operator_6_false_acc_9_nl));
  assign while_if_for_else_if_for_3_if_conc_1_pmx_7_4_lpi_2_dfm_1 = MUX_v_4_2_2(4'b0000,
      z_out_5, (z_out_8_7_2[5]));
  assign nl_operator_6_false_acc_10_nl = (operator_6_false_acc_2_cse_1[7:2]) + 6'b101111;
  assign operator_6_false_acc_10_nl = nl_operator_6_false_acc_10_nl[5:0];
  assign operator_6_false_acc_10_itm_5 = readslicef_6_1_5((operator_6_false_acc_10_nl));
  assign nl_operator_6_false_acc_8_nl = (operator_6_false_acc_2_cse_1[7:1]) + 7'b1011111;
  assign operator_6_false_acc_8_nl = nl_operator_6_false_acc_8_nl[6:0];
  assign operator_6_false_acc_8_itm_6_1 = readslicef_7_1_6((operator_6_false_acc_8_nl));
  assign nl_while_if_for_else_if_for_2_operator_6_false_acc_nl = conv_s2s_7_8({1'b1
      , (~ while_M_sva)}) + conv_u2s_7_8(while_if_for_t_7_0_sva_6_0);
  assign while_if_for_else_if_for_2_operator_6_false_acc_nl = nl_while_if_for_else_if_for_2_operator_6_false_acc_nl[7:0];
  assign while_if_for_else_if_for_2_operator_6_false_acc_itm_7_1 = readslicef_8_1_7((while_if_for_else_if_for_2_operator_6_false_acc_nl));
  assign nl_operator_6_false_acc_2_cse_1 = conv_u2u_7_8(while_if_for_t_7_0_sva_6_0)
      + conv_u2u_6_8(~ while_M_sva);
  assign operator_6_false_acc_2_cse_1 = nl_operator_6_false_acc_2_cse_1[7:0];
  assign nl_while_if_for_if_acc_nl = conv_u2s_4_5(while_if_for_t_7_0_sva_6_0[6:3])
      + 5'b11111;
  assign while_if_for_if_acc_nl = nl_while_if_for_if_acc_nl[4:0];
  assign while_if_for_if_acc_itm_4_1 = readslicef_5_1_4((while_if_for_if_acc_nl));
  assign while_if_for_asn_37 = ~(operator_6_false_slc_operator_6_false_acc_7_svs_mx1
      | while_if_for_if_acc_itm_4_1);
  assign while_if_for_asn_39 = operator_6_false_slc_operator_6_false_acc_7_svs_mx1
      & (~ while_if_for_if_acc_itm_4_1);
  assign or_tmp_7 = (fsm_output[4:3]!=2'b00);
  assign and_33_cse = (~ while_if_for_if_acc_itm_4_1) & (fsm_output[3]);
  assign and_37_cse = while_if_for_if_acc_itm_4_1 & (fsm_output[3]);
  assign while_if_for_if_for_if_while_if_for_if_for_if_and_cse = MUX_v_2_2_2(2'b00,
      (while_if_for_t_7_0_sva_6_0[4:3]), and_33_cse);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_psct_cse <= 1'b0;
      exit_while_if_for_sva <= 1'b0;
      while_if_for_t_7_0_sva_6_0 <= 7'b0000000;
      while_M_sva <= 6'b000000;
    end
    else if ( start_Pop_mioi_wen_comp ) begin
      reg_start_Pop_mioi_ccs_ccore_start_rsc_dat_ReadReqRun_psct_cse <= fsm_output[1];
      exit_while_if_for_sva <= ~ (readslicef_9_1_8((while_if_for_acc_nl)));
      while_if_for_t_7_0_sva_6_0 <= MUX_v_7_2_2(7'b0000000, (while_if_for_t_mux_1_nl),
          (not_nl));
      while_M_sva <= MUX_v_6_2_2(start_Pop_mioi_return_rsc_z, while_M_sva, or_tmp_7);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_6_false_slc_operator_6_false_acc_7_svs <= 1'b0;
    end
    else if ( start_Pop_mioi_wen_comp & (~(while_if_for_if_acc_itm_4_1 | (~ (fsm_output[3]))))
        ) begin
      operator_6_false_slc_operator_6_false_acc_7_svs <= operator_6_false_acc_itm_7_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      operator_33_true_return_6_0_sva <= 7'b0000000;
    end
    else if ( start_Pop_mioi_wen_comp & (~ or_tmp_7) ) begin
      operator_33_true_return_6_0_sva <= z_out_7[6:0];
    end
  end
  assign nl_while_if_for_acc_nl = conv_u2s_8_9(z_out_7) + conv_s2s_8_9({1'b1 , (~
      operator_33_true_return_6_0_sva)}) + 9'b000000001;
  assign while_if_for_acc_nl = nl_while_if_for_acc_nl[8:0];
  assign while_if_for_t_mux_1_nl = MUX_v_7_2_2((z_out_7[6:0]), while_if_for_t_7_0_sva_6_0,
      fsm_output[4]);
  assign not_nl = ~ (fsm_output[2]);
  assign while_if_for_if_for_if_mux_11_nl = MUX_v_3_2_2((while_if_for_t_7_0_sva_6_0[2:0]),
      (while_if_for_t_7_0_sva_6_0[4:2]), and_33_cse);
  assign nl_z_out = ({1'b1 , and_33_cse , 2'b11}) + conv_u2u_3_4(while_if_for_if_for_if_mux_11_nl);
  assign z_out = nl_z_out[3:0];
  assign while_if_for_else_if_for_if_mux_5_nl = MUX_v_4_2_2((while_if_for_t_7_0_sva_6_0[4:1]),
      (signext_4_3(while_if_for_t_7_0_sva_6_0[2:0])), and_37_cse);
  assign nl_z_out_1 = (while_if_for_else_if_for_if_mux_5_nl) + 4'b1101;
  assign z_out_1 = nl_z_out_1[3:0];
  assign not_42_nl = ~ and_33_cse;
  assign while_if_for_if_for_if_while_if_for_if_for_if_or_1_nl = MUX_v_2_2_2((while_if_for_t_7_0_sva_6_0[4:3]),
      2'b11, (not_42_nl));
  assign nl_z_out_2 = ({(while_if_for_if_for_if_while_if_for_if_for_if_or_1_nl) ,
      (while_if_for_t_7_0_sva_6_0[2:0])}) + conv_s2u_3_5({and_33_cse , 2'b01});
  assign z_out_2 = nl_z_out_2[4:0];
  assign nl_z_out_3 = ({while_if_for_if_for_if_while_if_for_if_for_if_and_cse , (while_if_for_t_7_0_sva_6_0[2:0])})
      + conv_s2u_4_5({1'b1 , (signext_2_1(~ and_33_cse)) , 1'b1});
  assign z_out_3 = nl_z_out_3[4:0];
  assign while_if_for_else_if_for_if_mux_6_nl = MUX_v_2_2_2((while_if_for_t_7_0_sva_6_0[4:3]),
      (signext_2_1(while_if_for_t_7_0_sva_6_0[2])), and_37_cse);
  assign nl_z_out_4 = ({(while_if_for_else_if_for_if_mux_6_nl) , (while_if_for_t_7_0_sva_6_0[2:0])})
      + conv_s2u_4_5({1'b1 , and_37_cse , 2'b11});
  assign z_out_4 = nl_z_out_4[4:0];
  assign nl_z_out_5 = ({while_if_for_if_for_if_while_if_for_if_for_if_and_cse , (while_if_for_t_7_0_sva_6_0[2:1])})
      + 4'b1111;
  assign z_out_5 = nl_z_out_5[3:0];
  assign nl_z_out_6 = ({while_if_for_if_for_if_while_if_for_if_for_if_and_cse , (while_if_for_t_7_0_sva_6_0[2:0])})
      + conv_s2u_3_5({1'b1 , and_33_cse , 1'b1});
  assign z_out_6 = nl_z_out_6[4:0];
  assign operator_6_false_mux_1_nl = MUX_v_7_2_2(({1'b0 , start_Pop_mioi_return_rsc_z}),
      while_if_for_t_7_0_sva_6_0, fsm_output[3]);
  assign nl_z_out_7 = conv_u2u_7_8(operator_6_false_mux_1_nl) + conv_u2u_3_8(signext_3_2({(fsm_output[2])
      , 1'b1}));
  assign z_out_7 = nl_z_out_7[7:0];
  assign while_if_for_if_for_if_mux_12_nl = MUX_v_8_2_2(({6'b111111 , (while_if_for_t_7_0_sva_6_0[2:1])}),
      operator_6_false_acc_2_cse_1, and_33_cse);
  assign nl_while_if_for_if_for_if_acc_nl = (while_if_for_if_for_if_mux_12_nl) +
      ({and_33_cse , 1'b0 , ({{4{and_33_cse}}, and_33_cse}) , 1'b1});
  assign while_if_for_if_for_if_acc_nl = nl_while_if_for_if_for_if_acc_nl[7:0];
  assign z_out_8_7_2 = readslicef_8_6_2((while_if_for_if_for_if_acc_nl));

  function automatic [0:0] MUX1HOT_s_1_3_2;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [2:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_3_2;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [2:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function automatic [3:0] MUX1HOT_v_4_3_2;
    input [3:0] input_2;
    input [3:0] input_1;
    input [3:0] input_0;
    input [2:0] sel;
    reg [3:0] result;
  begin
    result = input_0 & {4{sel[0]}};
    result = result | ( input_1 & {4{sel[1]}});
    result = result | ( input_2 & {4{sel[2]}});
    MUX1HOT_v_4_3_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [3:0] MUX_v_4_2_2;
    input [3:0] input_0;
    input [3:0] input_1;
    input [0:0] sel;
    reg [3:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_4_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [5:0] MUX_v_6_2_2;
    input [5:0] input_0;
    input [5:0] input_1;
    input [0:0] sel;
    reg [5:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_6_2_2 = result;
  end
  endfunction


  function automatic [6:0] MUX_v_7_2_2;
    input [6:0] input_0;
    input [6:0] input_1;
    input [0:0] sel;
    reg [6:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_7_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [0:0] readslicef_5_1_4;
    input [4:0] vector;
    reg [4:0] tmp;
  begin
    tmp = vector >> 4;
    readslicef_5_1_4 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_6_1_5;
    input [5:0] vector;
    reg [5:0] tmp;
  begin
    tmp = vector >> 5;
    readslicef_6_1_5 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_7_1_6;
    input [6:0] vector;
    reg [6:0] tmp;
  begin
    tmp = vector >> 6;
    readslicef_7_1_6 = tmp[0:0];
  end
  endfunction


  function automatic [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function automatic [5:0] readslicef_8_6_2;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 2;
    readslicef_8_6_2 = tmp[5:0];
  end
  endfunction


  function automatic [0:0] readslicef_9_1_8;
    input [8:0] vector;
    reg [8:0] tmp;
  begin
    tmp = vector >> 8;
    readslicef_9_1_8 = tmp[0:0];
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_2;
    input [1:0] vector;
  begin
    signext_3_2= {{1{vector[1]}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_1;
    input [0:0] vector;
  begin
    signext_4_1= {{3{vector[0]}}, vector};
  end
  endfunction


  function automatic [3:0] signext_4_3;
    input [2:0] vector;
  begin
    signext_4_3= {{1{vector[2]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_1;
    input [0:0] vector;
  begin
    signext_5_1= {{4{vector[0]}}, vector};
  end
  endfunction


  function automatic [4:0] signext_5_4;
    input [3:0] vector;
  begin
    signext_5_4= {{1{vector[3]}}, vector};
  end
  endfunction


  function automatic [7:0] conv_s2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_s2s_7_8 = {vector[6], vector};
  end
  endfunction


  function automatic [8:0] conv_s2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_s2s_8_9 = {vector[7], vector};
  end
  endfunction


  function automatic [4:0] conv_s2u_3_5 ;
    input [2:0]  vector ;
  begin
    conv_s2u_3_5 = {{2{vector[2]}}, vector};
  end
  endfunction


  function automatic [4:0] conv_s2u_4_5 ;
    input [3:0]  vector ;
  begin
    conv_s2u_4_5 = {vector[3], vector};
  end
  endfunction


  function automatic [4:0] conv_u2s_4_5 ;
    input [3:0]  vector ;
  begin
    conv_u2s_4_5 =  {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_8 =  {1'b0, vector};
  end
  endfunction


  function automatic [8:0] conv_u2s_8_9 ;
    input [7:0]  vector ;
  begin
    conv_u2s_8_9 =  {1'b0, vector};
  end
  endfunction


  function automatic [3:0] conv_u2u_3_4 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_4 = {1'b0, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_3_8 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_8 = {{5{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_6_8 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_8 = {{2{1'b0}}, vector};
  end
  endfunction


  function automatic [7:0] conv_u2u_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2u_7_8 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup_MemoryRun
// ------------------------------------------------------------------


module InputSetup_MemoryRun (
  clk, rst, write_req_val, write_req_rdy, write_req_msg, req_inter_val, req_inter_rdy,
      req_inter_msg, rsp_inter_val, rsp_inter_rdy, rsp_inter_msg, mem_inst_banks_bank_array_impl_data0_rsci_data_in_d,
      mem_inst_banks_bank_array_impl_data0_rsci_addr_d, mem_inst_banks_bank_array_impl_data0_rsci_re_d,
      mem_inst_banks_bank_array_impl_data0_rsci_we_d, mem_inst_banks_bank_array_impl_data0_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data0_rsci_en_d, mem_inst_banks_bank_array_impl_data1_rsci_data_in_d,
      mem_inst_banks_bank_array_impl_data1_rsci_addr_d, mem_inst_banks_bank_array_impl_data1_rsci_re_d,
      mem_inst_banks_bank_array_impl_data1_rsci_we_d, mem_inst_banks_bank_array_impl_data1_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data1_rsci_en_d, mem_inst_banks_bank_array_impl_data2_rsci_data_in_d,
      mem_inst_banks_bank_array_impl_data2_rsci_addr_d, mem_inst_banks_bank_array_impl_data2_rsci_re_d,
      mem_inst_banks_bank_array_impl_data2_rsci_we_d, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data2_rsci_en_d, mem_inst_banks_bank_array_impl_data3_rsci_data_in_d,
      mem_inst_banks_bank_array_impl_data3_rsci_addr_d, mem_inst_banks_bank_array_impl_data3_rsci_re_d,
      mem_inst_banks_bank_array_impl_data3_rsci_we_d, mem_inst_banks_bank_array_impl_data3_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data3_rsci_en_d, mem_inst_banks_bank_array_impl_data4_rsci_data_in_d,
      mem_inst_banks_bank_array_impl_data4_rsci_addr_d, mem_inst_banks_bank_array_impl_data4_rsci_re_d,
      mem_inst_banks_bank_array_impl_data4_rsci_we_d, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data4_rsci_en_d, mem_inst_banks_bank_array_impl_data5_rsci_data_in_d,
      mem_inst_banks_bank_array_impl_data5_rsci_addr_d, mem_inst_banks_bank_array_impl_data5_rsci_re_d,
      mem_inst_banks_bank_array_impl_data5_rsci_we_d, mem_inst_banks_bank_array_impl_data5_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data5_rsci_en_d, mem_inst_banks_bank_array_impl_data6_rsci_data_in_d,
      mem_inst_banks_bank_array_impl_data6_rsci_addr_d, mem_inst_banks_bank_array_impl_data6_rsci_re_d,
      mem_inst_banks_bank_array_impl_data6_rsci_we_d, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data6_rsci_en_d, mem_inst_banks_bank_array_impl_data7_rsci_data_in_d,
      mem_inst_banks_bank_array_impl_data7_rsci_addr_d, mem_inst_banks_bank_array_impl_data7_rsci_re_d,
      mem_inst_banks_bank_array_impl_data7_rsci_we_d, mem_inst_banks_bank_array_impl_data7_rsci_data_out_d,
      mem_inst_banks_bank_array_impl_data7_rsci_en_d
);
  input clk;
  input rst;
  input write_req_val;
  output write_req_rdy;
  input [68:0] write_req_msg;
  input req_inter_val;
  output req_inter_rdy;
  input [136:0] req_inter_msg;
  output rsp_inter_val;
  input rsp_inter_rdy;
  output [71:0] rsp_inter_msg;
  output [7:0] mem_inst_banks_bank_array_impl_data0_rsci_data_in_d;
  output [4:0] mem_inst_banks_bank_array_impl_data0_rsci_addr_d;
  output mem_inst_banks_bank_array_impl_data0_rsci_re_d;
  output mem_inst_banks_bank_array_impl_data0_rsci_we_d;
  input [7:0] mem_inst_banks_bank_array_impl_data0_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data0_rsci_en_d;
  output [7:0] mem_inst_banks_bank_array_impl_data1_rsci_data_in_d;
  output [4:0] mem_inst_banks_bank_array_impl_data1_rsci_addr_d;
  output mem_inst_banks_bank_array_impl_data1_rsci_re_d;
  output mem_inst_banks_bank_array_impl_data1_rsci_we_d;
  input [7:0] mem_inst_banks_bank_array_impl_data1_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data1_rsci_en_d;
  output [7:0] mem_inst_banks_bank_array_impl_data2_rsci_data_in_d;
  output [4:0] mem_inst_banks_bank_array_impl_data2_rsci_addr_d;
  output mem_inst_banks_bank_array_impl_data2_rsci_re_d;
  output mem_inst_banks_bank_array_impl_data2_rsci_we_d;
  input [7:0] mem_inst_banks_bank_array_impl_data2_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data2_rsci_en_d;
  output [7:0] mem_inst_banks_bank_array_impl_data3_rsci_data_in_d;
  output [4:0] mem_inst_banks_bank_array_impl_data3_rsci_addr_d;
  output mem_inst_banks_bank_array_impl_data3_rsci_re_d;
  output mem_inst_banks_bank_array_impl_data3_rsci_we_d;
  input [7:0] mem_inst_banks_bank_array_impl_data3_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data3_rsci_en_d;
  output [7:0] mem_inst_banks_bank_array_impl_data4_rsci_data_in_d;
  output [4:0] mem_inst_banks_bank_array_impl_data4_rsci_addr_d;
  output mem_inst_banks_bank_array_impl_data4_rsci_re_d;
  output mem_inst_banks_bank_array_impl_data4_rsci_we_d;
  input [7:0] mem_inst_banks_bank_array_impl_data4_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data4_rsci_en_d;
  output [7:0] mem_inst_banks_bank_array_impl_data5_rsci_data_in_d;
  output [4:0] mem_inst_banks_bank_array_impl_data5_rsci_addr_d;
  output mem_inst_banks_bank_array_impl_data5_rsci_re_d;
  output mem_inst_banks_bank_array_impl_data5_rsci_we_d;
  input [7:0] mem_inst_banks_bank_array_impl_data5_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data5_rsci_en_d;
  output [7:0] mem_inst_banks_bank_array_impl_data6_rsci_data_in_d;
  output [4:0] mem_inst_banks_bank_array_impl_data6_rsci_addr_d;
  output mem_inst_banks_bank_array_impl_data6_rsci_re_d;
  output mem_inst_banks_bank_array_impl_data6_rsci_we_d;
  input [7:0] mem_inst_banks_bank_array_impl_data6_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data6_rsci_en_d;
  output [7:0] mem_inst_banks_bank_array_impl_data7_rsci_data_in_d;
  output [4:0] mem_inst_banks_bank_array_impl_data7_rsci_addr_d;
  output mem_inst_banks_bank_array_impl_data7_rsci_re_d;
  output mem_inst_banks_bank_array_impl_data7_rsci_we_d;
  input [7:0] mem_inst_banks_bank_array_impl_data7_rsci_data_out_d;
  output mem_inst_banks_bank_array_impl_data7_rsci_en_d;


  // Interconnect Declarations
  wire MemoryRun_wten;
  wire req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt;
  wire [7:0] req_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
  wire [63:0] req_inter_PopNB_mioi_data_addr_rsc_z_mxwt;
  wire [63:0] req_inter_PopNB_mioi_data_data_rsc_z_mxwt;
  wire req_inter_PopNB_mioi_return_rsc_z_mxwt;
  wire [63:0] write_req_PopNB_mioi_data_data_data_rsc_z_mxwt;
  wire [4:0] write_req_PopNB_mioi_data_index_rsc_z_mxwt;
  wire write_req_PopNB_mioi_return_rsc_z_mxwt;
  wire rsp_inter_Push_mioi_wen_comp;
  wire [7:0] mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg;
  wire [7:0] mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg;
  wire [7:0] mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg;
  wire [7:0] mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg;
  wire [7:0] mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg;
  wire [7:0] mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg;
  wire [7:0] mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg;
  wire [7:0] mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg;
  wire [1:0] fsm_output;
  wire mem_inst_request_xbar_xbar_for_3_if_1_mux_28_tmp;
  wire mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp;
  wire mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp;
  wire mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp;
  wire mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp;
  wire mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp;
  wire mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp;
  wire mem_inst_request_xbar_xbar_for_3_if_1_mux_tmp;
  wire [7:0] mem_inst_request_xbar_xbar_for_8_lshift_tmp;
  wire [7:0] mem_inst_request_xbar_xbar_for_7_lshift_tmp;
  wire [7:0] mem_inst_request_xbar_xbar_for_6_lshift_tmp;
  wire [7:0] mem_inst_request_xbar_xbar_for_5_lshift_tmp;
  wire [7:0] mem_inst_request_xbar_xbar_for_4_lshift_tmp;
  wire [7:0] mem_inst_request_xbar_xbar_for_3_lshift_tmp;
  wire [7:0] mem_inst_request_xbar_xbar_for_2_lshift_tmp;
  wire [7:0] mem_inst_request_xbar_xbar_for_1_lshift_tmp;
  wire while_if_1_while_if_1_or_tmp;
  wire and_dcpl;
  wire and_dcpl_1;
  wire or_dcpl_1;
  wire nor_tmp_1;
  wire and_tmp;
  wire and_tmp_1;
  wire and_tmp_2;
  wire and_tmp_3;
  wire and_tmp_4;
  wire and_tmp_5;
  wire and_tmp_6;
  wire and_tmp_7;
  wire or_dcpl_11;
  wire or_dcpl_12;
  wire and_dcpl_122;
  wire and_dcpl_131;
  wire and_dcpl_134;
  wire and_dcpl_144;
  wire and_dcpl_148;
  wire and_dcpl_151;
  wire and_dcpl_157;
  wire and_dcpl_167;
  wire and_dcpl_171;
  wire or_dcpl_24;
  wire or_dcpl_27;
  wire or_dcpl_30;
  wire or_dcpl_33;
  wire or_dcpl_36;
  wire or_dcpl_39;
  wire or_dcpl_40;
  wire or_dcpl_41;
  wire or_dcpl_42;
  wire or_dcpl_43;
  wire or_dcpl_44;
  wire or_dcpl_45;
  wire or_dcpl_47;
  wire and_dcpl_185;
  wire or_dcpl_49;
  wire or_dcpl_50;
  wire or_dcpl_51;
  wire or_dcpl_52;
  wire and_dcpl_189;
  wire and_dcpl_190;
  wire or_dcpl_53;
  wire or_dcpl_54;
  wire or_dcpl_55;
  wire or_dcpl_56;
  wire or_dcpl_57;
  wire and_dcpl_206;
  wire or_dcpl_61;
  wire or_dcpl_62;
  wire or_dcpl_63;
  wire or_dcpl_64;
  wire and_dcpl_210;
  wire and_dcpl_213;
  wire or_dcpl_65;
  wire or_dcpl_66;
  wire or_dcpl_67;
  wire or_dcpl_68;
  wire or_dcpl_69;
  wire and_dcpl_229;
  wire or_dcpl_73;
  wire or_dcpl_74;
  wire or_dcpl_75;
  wire or_dcpl_76;
  wire and_dcpl_233;
  wire and_dcpl_236;
  wire or_dcpl_77;
  wire or_dcpl_78;
  wire or_dcpl_79;
  wire or_dcpl_80;
  wire or_dcpl_81;
  wire and_dcpl_252;
  wire or_dcpl_85;
  wire or_dcpl_86;
  wire or_dcpl_87;
  wire or_dcpl_88;
  wire and_dcpl_256;
  wire and_dcpl_259;
  wire or_dcpl_89;
  wire or_dcpl_90;
  wire or_dcpl_91;
  wire or_dcpl_92;
  wire or_dcpl_93;
  wire and_dcpl_275;
  wire or_dcpl_97;
  wire or_dcpl_98;
  wire or_dcpl_99;
  wire or_dcpl_100;
  wire and_dcpl_279;
  wire and_dcpl_281;
  wire or_dcpl_101;
  wire or_dcpl_102;
  wire or_dcpl_103;
  wire or_dcpl_104;
  wire or_dcpl_105;
  wire or_dcpl_107;
  wire and_dcpl_297;
  wire or_dcpl_109;
  wire or_dcpl_110;
  wire or_dcpl_111;
  wire or_dcpl_112;
  wire and_dcpl_301;
  wire and_dcpl_302;
  wire or_dcpl_113;
  wire or_dcpl_114;
  wire or_dcpl_115;
  wire or_dcpl_116;
  wire or_dcpl_117;
  wire and_dcpl_318;
  wire or_dcpl_121;
  wire or_dcpl_122;
  wire or_dcpl_123;
  wire or_dcpl_124;
  wire and_dcpl_322;
  wire and_dcpl_323;
  wire or_dcpl_125;
  wire or_dcpl_126;
  wire or_dcpl_127;
  wire or_dcpl_128;
  wire or_dcpl_129;
  wire or_dcpl_131;
  wire and_dcpl_339;
  wire or_dcpl_133;
  wire or_dcpl_134;
  wire or_dcpl_135;
  wire or_dcpl_136;
  wire and_dcpl_343;
  wire and_dcpl_344;
  wire or_dcpl_137;
  wire mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
  wire Arbiter_8U_Roundrobin_pick_unequal_tmp_15;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_lpi_1_dfm_mx0;
  wire operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_11_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_10_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_14_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_13_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_12_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_9_sva_1;
  reg mem_inst_request_xbar_arbiters_next_7_1_sva;
  reg mem_inst_request_xbar_arbiters_next_7_3_sva;
  reg mem_inst_request_xbar_arbiters_next_7_4_sva;
  reg mem_inst_request_xbar_arbiters_next_7_2_sva;
  reg mem_inst_request_xbar_arbiters_next_7_5_sva;
  reg mem_inst_request_xbar_arbiters_next_7_6_sva;
  reg mem_inst_request_xbar_arbiters_next_7_7_sva;
  wire Arbiter_8U_Roundrobin_pick_unequal_tmp_14;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_7_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_7_lpi_1_dfm_mx0;
  wire operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_11_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_10_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_14_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_13_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_12_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_9_7_sva_1;
  reg mem_inst_request_xbar_arbiters_next_6_1_sva;
  reg mem_inst_request_xbar_arbiters_next_6_3_sva;
  reg mem_inst_request_xbar_arbiters_next_6_4_sva;
  reg mem_inst_request_xbar_arbiters_next_6_2_sva;
  reg mem_inst_request_xbar_arbiters_next_6_5_sva;
  reg mem_inst_request_xbar_arbiters_next_6_6_sva;
  reg mem_inst_request_xbar_arbiters_next_6_7_sva;
  wire Arbiter_8U_Roundrobin_pick_unequal_tmp_13;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_6_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_6_lpi_1_dfm_mx0;
  wire operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_11_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_10_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_13_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_12_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_9_6_sva_1;
  reg mem_inst_request_xbar_arbiters_next_5_1_sva;
  reg mem_inst_request_xbar_arbiters_next_5_3_sva;
  reg mem_inst_request_xbar_arbiters_next_5_4_sva;
  reg mem_inst_request_xbar_arbiters_next_5_2_sva;
  reg mem_inst_request_xbar_arbiters_next_5_5_sva;
  reg mem_inst_request_xbar_arbiters_next_5_6_sva;
  reg mem_inst_request_xbar_arbiters_next_5_7_sva;
  wire Arbiter_8U_Roundrobin_pick_unequal_tmp_12;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_5_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_5_lpi_1_dfm_mx0;
  wire operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_11_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_10_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_14_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_13_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_12_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_9_5_sva_1;
  reg mem_inst_request_xbar_arbiters_next_4_1_sva;
  reg mem_inst_request_xbar_arbiters_next_4_3_sva;
  reg mem_inst_request_xbar_arbiters_next_4_4_sva;
  reg mem_inst_request_xbar_arbiters_next_4_2_sva;
  reg mem_inst_request_xbar_arbiters_next_4_5_sva;
  reg mem_inst_request_xbar_arbiters_next_4_6_sva;
  reg mem_inst_request_xbar_arbiters_next_4_7_sva;
  wire Arbiter_8U_Roundrobin_pick_unequal_tmp_11;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_4_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_4_lpi_1_dfm_mx0;
  wire operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_11_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_10_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_14_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_13_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_12_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_9_4_sva_1;
  reg mem_inst_request_xbar_arbiters_next_3_1_sva;
  reg mem_inst_request_xbar_arbiters_next_3_3_sva;
  reg mem_inst_request_xbar_arbiters_next_3_4_sva;
  reg mem_inst_request_xbar_arbiters_next_3_2_sva;
  reg mem_inst_request_xbar_arbiters_next_3_5_sva;
  reg mem_inst_request_xbar_arbiters_next_3_6_sva;
  reg mem_inst_request_xbar_arbiters_next_3_7_sva;
  wire Arbiter_8U_Roundrobin_pick_unequal_tmp_10;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_3_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_3_lpi_1_dfm_mx0;
  wire operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_11_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_10_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_14_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_13_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_12_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_9_3_sva_1;
  reg mem_inst_request_xbar_arbiters_next_2_1_sva;
  reg mem_inst_request_xbar_arbiters_next_2_3_sva;
  reg mem_inst_request_xbar_arbiters_next_2_4_sva;
  reg mem_inst_request_xbar_arbiters_next_2_2_sva;
  reg mem_inst_request_xbar_arbiters_next_2_5_sva;
  reg mem_inst_request_xbar_arbiters_next_2_6_sva;
  reg mem_inst_request_xbar_arbiters_next_2_7_sva;
  wire Arbiter_8U_Roundrobin_pick_unequal_tmp_9;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_2_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_2_lpi_1_dfm_mx0;
  wire operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_11_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_10_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_14_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_13_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_12_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_9_2_sva_1;
  reg mem_inst_request_xbar_arbiters_next_1_1_sva;
  reg mem_inst_request_xbar_arbiters_next_1_3_sva;
  reg mem_inst_request_xbar_arbiters_next_1_4_sva;
  reg mem_inst_request_xbar_arbiters_next_1_2_sva;
  reg mem_inst_request_xbar_arbiters_next_1_5_sva;
  reg mem_inst_request_xbar_arbiters_next_1_6_sva;
  reg mem_inst_request_xbar_arbiters_next_1_7_sva;
  wire Arbiter_8U_Roundrobin_pick_unequal_tmp_8;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_1_lpi_1_dfm_mx0;
  wire nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_1_lpi_1_dfm_mx0;
  wire operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_11_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_10_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_14_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_13_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_12_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_priority_9_1_sva_1;
  reg mem_inst_request_xbar_arbiters_next_0_1_sva;
  reg mem_inst_request_xbar_arbiters_next_0_3_sva;
  reg mem_inst_request_xbar_arbiters_next_0_4_sva;
  reg mem_inst_request_xbar_arbiters_next_0_2_sva;
  reg mem_inst_request_xbar_arbiters_next_0_5_sva;
  reg mem_inst_request_xbar_arbiters_next_0_6_sva;
  reg mem_inst_request_xbar_arbiters_next_0_7_sva;
  reg while_asn_mdf_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1;
  wire mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  wire mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  wire mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  wire mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  wire mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  wire mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  wire mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1;
  wire [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_1;
  wire mem_inst_load_store_valid_src_7_lpi_1_dfm_7_mx0;
  wire [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_1;
  wire mem_inst_load_store_valid_src_6_lpi_1_dfm_7_mx0;
  wire [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_1;
  wire mem_inst_load_store_valid_src_5_lpi_1_dfm_7_mx0;
  wire [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_1;
  wire mem_inst_load_store_valid_src_4_lpi_1_dfm_7_mx0;
  wire [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_1;
  wire mem_inst_load_store_valid_src_3_lpi_1_dfm_7_mx0;
  wire [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_1;
  wire mem_inst_load_store_valid_src_2_lpi_1_dfm_7_mx0;
  wire [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_1;
  wire mem_inst_load_store_valid_src_1_lpi_1_dfm_7_mx0;
  wire [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_1;
  wire mem_inst_load_store_valid_src_0_lpi_1_dfm_7_mx0;
  wire mem_inst_load_store_valid_src_7_lpi_1_dfm_8;
  wire mem_inst_load_store_for_4_if_and_tmp_8_sva_1;
  wire mem_inst_load_store_valid_src_6_lpi_1_dfm_8;
  wire mem_inst_load_store_for_4_if_and_tmp_9_sva_1;
  wire mem_inst_load_store_valid_src_5_lpi_1_dfm_8;
  wire mem_inst_load_store_for_4_if_and_tmp_10_sva_1;
  wire mem_inst_load_store_valid_src_4_lpi_1_dfm_8;
  wire mem_inst_load_store_for_4_if_and_tmp_11_sva_1;
  wire mem_inst_load_store_valid_src_3_lpi_1_dfm_8;
  wire mem_inst_load_store_for_4_if_and_tmp_12_sva_1;
  wire mem_inst_load_store_valid_src_2_lpi_1_dfm_8;
  wire mem_inst_load_store_for_4_if_and_tmp_13_sva_1;
  wire mem_inst_load_store_valid_src_1_lpi_1_dfm_8;
  wire mem_inst_load_store_for_4_if_and_tmp_14_sva_1;
  wire mem_inst_load_store_valid_src_0_lpi_1_dfm_8;
  wire mem_inst_load_store_for_4_if_and_tmp_15_sva_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_7_sva_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_7_sva_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_7_sva_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_7_sva_1;
  wire mem_inst_load_store_for_4_if_and_tmp_sva_2;
  wire mem_inst_load_store_for_4_and_55_cse_1;
  wire mem_inst_load_store_for_4_and_7_tmp_1;
  wire mem_inst_load_store_for_4_and_15_tmp_1;
  wire mem_inst_load_store_for_4_and_23_tmp_1;
  wire mem_inst_load_store_for_4_and_31_tmp_1;
  wire mem_inst_load_store_for_4_and_39_tmp_1;
  wire mem_inst_load_store_for_4_if_and_tmp_1_sva_2;
  wire mem_inst_load_store_for_4_and_53_cse_1;
  wire mem_inst_load_store_for_4_and_6_tmp_1;
  wire mem_inst_load_store_for_4_and_14_tmp_1;
  wire mem_inst_load_store_for_4_and_22_tmp_1;
  wire mem_inst_load_store_for_4_and_30_tmp_1;
  wire mem_inst_load_store_for_4_and_38_tmp_1;
  wire mem_inst_load_store_for_4_if_and_tmp_2_sva_2;
  wire mem_inst_load_store_for_4_and_51_cse_1;
  wire mem_inst_load_store_for_4_and_5_tmp_1;
  wire mem_inst_load_store_for_4_and_13_tmp_1;
  wire mem_inst_load_store_for_4_and_21_tmp_1;
  wire mem_inst_load_store_for_4_and_29_tmp_1;
  wire mem_inst_load_store_for_4_and_37_tmp_1;
  wire mem_inst_load_store_for_4_if_and_tmp_3_sva_2;
  wire mem_inst_load_store_for_4_and_49_cse_1;
  wire mem_inst_load_store_for_4_and_4_tmp_1;
  wire mem_inst_load_store_for_4_and_12_tmp_1;
  wire mem_inst_load_store_for_4_and_20_tmp_1;
  wire mem_inst_load_store_for_4_and_28_tmp_1;
  wire mem_inst_load_store_for_4_and_36_tmp_1;
  wire mem_inst_load_store_for_4_if_and_tmp_4_sva_2;
  wire mem_inst_load_store_for_4_and_47_cse_1;
  wire mem_inst_load_store_for_4_and_3_tmp_1;
  wire mem_inst_load_store_for_4_and_11_tmp_1;
  wire mem_inst_load_store_for_4_and_19_tmp_1;
  wire mem_inst_load_store_for_4_and_27_tmp_1;
  wire mem_inst_load_store_for_4_and_35_tmp_1;
  wire mem_inst_load_store_for_4_if_and_tmp_5_sva_2;
  wire mem_inst_load_store_for_4_and_45_cse_1;
  wire mem_inst_load_store_for_4_and_2_tmp_1;
  wire mem_inst_load_store_for_4_and_10_tmp_1;
  wire mem_inst_load_store_for_4_and_18_tmp_1;
  wire mem_inst_load_store_for_4_and_26_tmp_1;
  wire mem_inst_load_store_for_4_and_34_tmp_1;
  wire mem_inst_load_store_for_4_if_and_tmp_6_sva_2;
  wire mem_inst_load_store_for_4_and_43_cse_1;
  wire mem_inst_load_store_for_4_and_1_tmp_1;
  wire mem_inst_load_store_for_4_and_9_tmp_1;
  wire mem_inst_load_store_for_4_and_17_tmp_1;
  wire mem_inst_load_store_for_4_and_25_tmp_1;
  wire mem_inst_load_store_for_4_and_33_tmp_1;
  wire mem_inst_load_store_for_4_if_and_tmp_7_sva_2;
  wire mem_inst_load_store_for_4_and_41_cse_1;
  wire mem_inst_load_store_for_4_and_tmp_1;
  wire mem_inst_load_store_for_4_and_8_tmp_1;
  wire mem_inst_load_store_for_4_and_16_tmp_1;
  wire mem_inst_load_store_for_4_and_24_tmp_1;
  wire mem_inst_load_store_for_4_and_32_tmp_1;
  wire mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_23_m1c_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_1_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_6_sva_mx1;
  wire mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_22_m1c_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_1_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_6_sva_mx1;
  wire mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_21_m1c_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_1_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_6_sva_mx1;
  wire mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_20_m1c_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_1_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_6_sva_mx1;
  wire mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_19_m1c_1;
  wire mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_18_m1c_1;
  wire mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_17_m1c_1;
  wire mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_16_m1c_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_4_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_5_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_4_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_5_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_4_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_5_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_4_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_5_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_2_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_3_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_2_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_3_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_2_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_3_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_2_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_3_sva_mx1;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_sva_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_sva_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_sva_1;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_sva_1;
  reg while_stage_0_3;
  reg while_asn_mdf_sva_st_1_2;
  reg while_lor_lpi_1_dfm_st_1;
  reg while_lor_lpi_1_dfm_2;
  reg mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1;
  reg mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1;
  reg mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1;
  reg mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1;
  reg mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1;
  reg mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1;
  reg mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1;
  reg mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1;
  reg while_stage_0_5;
  wire one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_sva_1;
  wire one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_sva_1;
  wire one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_sva_1;
  wire one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_7_sva_1;
  wire one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_7_sva_1;
  wire one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_7_sva_1;
  wire one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_6_sva_1;
  wire one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_6_sva_1;
  wire one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_6_sva_1;
  wire one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_5_sva_1;
  wire one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_5_sva_1;
  wire one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_5_sva_1;
  wire one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_4_sva_1;
  wire one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_4_sva_1;
  wire one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_4_sva_1;
  wire one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_3_sva_1;
  wire one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_3_sva_1;
  wire one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_3_sva_1;
  wire one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_2_sva_1;
  wire one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_2_sva_1;
  wire one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_2_sva_1;
  wire one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_1_sva_1;
  wire one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_1_sva_1;
  wire one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_1_sva_1;
  wire [2:0] mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2;
  wire mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2;
  wire mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2;
  wire mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2;
  wire mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2;
  wire mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2;
  wire mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2;
  wire [2:0] mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1;
  wire [2:0] mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx0w0;
  wire [2:0] mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx0w0;
  wire [2:0] mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx0w0;
  wire [2:0] mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx0w0;
  wire [2:0] mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx0w0;
  wire [2:0] mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx0w0;
  reg reg_mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_ftd;
  reg reg_mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_ftd;
  reg reg_mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_ftd;
  reg reg_mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_ftd;
  reg reg_mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_ftd;
  reg reg_mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_ftd;
  wire mem_inst_banks_read_for_mux_cse;
  wire mem_inst_banks_write_if_for_if_mux_cse;
  wire mem_inst_banks_read_for_mux_4_cse;
  wire mem_inst_banks_write_if_for_if_mux_4_cse;
  wire mem_inst_banks_read_for_mux_8_cse;
  wire mem_inst_banks_write_if_for_if_mux_8_cse;
  wire mem_inst_banks_read_for_mux_12_cse;
  wire mem_inst_banks_write_if_for_if_mux_12_cse;
  wire mem_inst_banks_read_for_mux_16_cse;
  wire mem_inst_banks_write_if_for_if_mux_16_cse;
  wire mem_inst_banks_read_for_mux_20_cse;
  wire mem_inst_banks_write_if_for_if_mux_20_cse;
  wire mem_inst_banks_read_for_mux_24_cse;
  wire mem_inst_banks_write_if_for_if_mux_24_cse;
  wire mem_inst_banks_read_for_mux_28_cse;
  wire mem_inst_banks_write_if_for_if_mux_28_cse;
  reg reg_rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse;
  reg reg_write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse;
  reg reg_req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse;
  reg reg_mem_inst_banks_bank_array_impl_data7_rsc_cgo_cse;
  reg reg_mem_inst_banks_bank_array_impl_data6_rsc_cgo_cse;
  reg reg_mem_inst_banks_bank_array_impl_data5_rsc_cgo_cse;
  reg reg_mem_inst_banks_bank_array_impl_data4_rsc_cgo_cse;
  reg reg_mem_inst_banks_bank_array_impl_data3_rsc_cgo_cse;
  reg reg_mem_inst_banks_bank_array_impl_data2_rsc_cgo_cse;
  reg reg_mem_inst_banks_bank_array_impl_data1_rsc_cgo_cse;
  reg reg_mem_inst_banks_bank_array_impl_data0_rsc_cgo_cse;
  wire mem_inst_request_xbar_arbiters_next_and_cse;
  wire mem_inst_request_xbar_arbiters_next_and_7_cse;
  wire mem_inst_request_xbar_arbiters_next_and_14_cse;
  wire mem_inst_request_xbar_arbiters_next_and_21_cse;
  wire mem_inst_request_xbar_arbiters_next_and_28_cse;
  wire mem_inst_request_xbar_arbiters_next_and_35_cse;
  wire mem_inst_request_xbar_arbiters_next_and_42_cse;
  wire operator_15_false_and_cse;
  wire crossbar_InputSetup_InputType_8U_8U_for_aelse_and_cse;
  wire mem_inst_load_store_for_4_if_and_104_cse;
  wire mem_inst_load_store_for_4_if_and_108_cse;
  wire mem_inst_load_store_for_4_if_and_112_cse;
  wire mem_inst_load_store_for_4_if_and_116_cse;
  wire mem_inst_load_store_for_4_if_and_120_cse;
  wire mem_inst_load_store_for_4_if_and_124_cse;
  wire and_685_cse;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1;
  wire and_525_rmff;
  wire and_523_rmff;
  wire and_521_rmff;
  wire and_519_rmff;
  wire and_517_rmff;
  wire and_515_rmff;
  wire and_513_rmff;
  wire and_511_rmff;
  wire MemoryRun_wten_iff;
  wire and_231_rmff;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1_dfm_1_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1_dfm_1_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1_dfm_1_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1_dfm_1_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1_dfm_1_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1_dfm_1_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1_dfm_1_2;
  reg [7:0] crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1;
  wire [7:0] crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2;
  reg [7:0] crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1;
  wire [7:0] crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2;
  reg [7:0] crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1;
  wire [7:0] crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2;
  reg [7:0] crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1;
  wire [7:0] crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2;
  reg [7:0] crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1;
  wire [7:0] crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2;
  reg [7:0] crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1;
  wire [7:0] crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2;
  reg [7:0] crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1;
  wire [7:0] crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2;
  reg [7:0] mem_inst_load_store_data_out_0_lpi_1_dfm_1;
  wire [7:0] mem_inst_load_store_data_out_0_lpi_1_dfm_2;
  wire [7:0] while_req_reg_data_0_lpi_1_dfm_1_mx0;
  wire [7:0] while_req_reg_data_1_lpi_1_dfm_1_mx0;
  wire [7:0] while_req_reg_data_2_lpi_1_dfm_1_mx0;
  wire [7:0] while_req_reg_data_3_lpi_1_dfm_1_mx0;
  wire [7:0] while_req_reg_data_4_lpi_1_dfm_1_mx0;
  wire [7:0] while_req_reg_data_5_lpi_1_dfm_1_mx0;
  wire [7:0] while_req_reg_data_6_lpi_1_dfm_1_mx0;
  wire [7:0] while_req_reg_data_7_lpi_1_dfm_1_mx0;
  wire [4:0] while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0;
  wire [4:0] while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0;
  wire [4:0] while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0;
  wire [4:0] while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0;
  wire [4:0] while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0;
  wire [4:0] while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0;
  wire [4:0] while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0;
  wire [4:0] while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0;
  reg [63:0] while_req_reg_addr_sva_1;
  wire and_687_tmp;
  wire and_688_tmp;
  wire and_689_tmp;
  wire and_690_tmp;
  wire and_691_tmp;
  wire and_692_tmp;
  wire and_693_tmp;
  wire and_694_tmp;
  wire while_and_itm;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_3;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_4;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_5;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_6;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_7;
  wire Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_7;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1;
  reg mem_inst_load_store_for_4_if_and_stg_1_3_1_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_2_1_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_1_1_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_0_1_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_3_2_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_2_2_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_1_2_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_0_2_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_3_3_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_2_3_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_1_3_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_0_3_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_3_4_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_2_4_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_1_4_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_0_4_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_3_5_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_2_5_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_1_5_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_0_5_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_3_6_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_2_6_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_1_6_sva;
  reg mem_inst_load_store_for_4_if_and_stg_1_0_6_sva;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1;
  reg while_stage_0_4;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1_dfm_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1_dfm_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1_dfm_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1_dfm_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1_dfm_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1_dfm_2;
  reg crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1_dfm_2;
  reg while_req_reg_type_val_sva_1;
  reg [7:0] while_req_reg_valids_sva_1;
  reg [63:0] while_req_reg_data_sva_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_2;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_1_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_2;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_1_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_2;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_1_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_2;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_1_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_2;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_1_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_2;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_1_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_2;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_1_1;
  reg [2:0] crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_2;
  reg while_asn_mdf_sva_st_1_3;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_1_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_1_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_1_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_1_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_2_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_2_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_2_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_2_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_3_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_3_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_3_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_3_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_4_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_4_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_4_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_4_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_5_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_5_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_5_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_5_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_0_6_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_1_6_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_2_6_sva_mx0w0;
  wire mem_inst_load_store_for_4_if_and_stg_1_3_6_sva_mx0w0;
  wire mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1;
  wire mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1;
  wire mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1;
  wire mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1;
  wire mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1;
  wire mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1;
  wire mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1;
  wire mem_inst_compute_bank_request_for_land_lpi_1_dfm_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1;
  wire mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
  wire operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1;
  wire operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1;
  wire operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1;
  wire while_req_reg_valids_7_lpi_1_dfm_1_mx0;
  wire while_req_reg_valids_6_lpi_1_dfm_1_mx0;
  wire while_and_21_cse_1;
  wire while_req_reg_valids_5_lpi_1_dfm_1_mx0;
  wire while_req_reg_valids_4_lpi_1_dfm_1_mx0;
  wire while_req_reg_valids_3_lpi_1_dfm_1_mx0;
  wire while_req_reg_valids_2_lpi_1_dfm_1_mx0;
  wire while_req_reg_valids_1_lpi_1_dfm_1_mx0;
  wire while_req_reg_valids_0_lpi_1_dfm_1_mx0;
  wire while_req_reg_type_val_lpi_1_dfm_2;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1;
  wire Arbiter_8U_Roundrobin_pick_if_1_not_64;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1;
  wire mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0;
  wire crossbar_InputSetup_InputType_8U_8U_for_aelse_and_8_cse;
  wire crossbar_InputSetup_InputType_8U_8U_for_and_7_cse;
  wire crossbar_InputSetup_InputType_8U_8U_for_aelse_and_16_cse;
  wire mem_inst_request_xbar_xbar_for_3_and_cse;
  wire while_req_reg_addr_and_cse;
  wire while_oelse_and_1_cse;
  wire crossbar_InputSetup_InputType_8U_8U_for_and_20_cse;

  wire[0:0] and_30_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb;
  wire[0:0] and_32_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1;
  wire[0:0] and_35_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2;
  wire[0:0] and_37_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3;
  wire[0:0] and_40_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4;
  wire[0:0] and_42_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5;
  wire[0:0] and_45_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6;
  wire[0:0] and_47_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7;
  wire[0:0] and_50_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8;
  wire[0:0] and_52_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9;
  wire[0:0] and_55_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10;
  wire[0:0] and_57_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11;
  wire[0:0] and_60_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12;
  wire[0:0] and_62_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13;
  wire[0:0] and_65_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14;
  wire[0:0] and_67_nl;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15;
  wire[0:0] pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15;
  wire[0:0] pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15;
  wire[0:0] mux_nl;
  wire[0:0] or_2_nl;
  wire[0:0] crossbar_InputSetup_InputType_8U_8U_for_mux_27_nl;
  wire[0:0] crossbar_InputSetup_InputType_8U_8U_for_mux_25_nl;
  wire[0:0] crossbar_InputSetup_InputType_8U_8U_for_mux_23_nl;
  wire[0:0] crossbar_InputSetup_InputType_8U_8U_for_mux_21_nl;
  wire[0:0] crossbar_InputSetup_InputType_8U_8U_for_mux_19_nl;
  wire[0:0] crossbar_InputSetup_InputType_8U_8U_for_mux_17_nl;
  wire[0:0] crossbar_InputSetup_InputType_8U_8U_for_mux_14_nl;
  wire[0:0] crossbar_InputSetup_InputType_8U_8U_for_mux_29_nl;
  wire[2:0] crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_14_nl;
  wire[1:0] mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_7_nl;
  wire[0:0] mem_inst_load_store_for_4_and_116_nl;
  wire[0:0] mem_inst_load_store_for_4_and_71_nl;
  wire[0:0] mem_inst_load_store_for_4_and_117_nl;
  wire[0:0] mem_inst_load_store_for_4_and_87_nl;
  wire[0:0] mem_inst_load_store_for_4_and_102_nl;
  wire[0:0] and_695_nl;
  wire[2:0] crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_12_nl;
  wire[1:0] mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_6_nl;
  wire[0:0] mem_inst_load_store_for_4_and_114_nl;
  wire[0:0] mem_inst_load_store_for_4_and_69_nl;
  wire[0:0] mem_inst_load_store_for_4_and_115_nl;
  wire[0:0] mem_inst_load_store_for_4_and_85_nl;
  wire[0:0] mem_inst_load_store_for_4_and_100_nl;
  wire[0:0] and_696_nl;
  wire[2:0] crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_10_nl;
  wire[1:0] mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_5_nl;
  wire[0:0] mem_inst_load_store_for_4_and_112_nl;
  wire[0:0] mem_inst_load_store_for_4_and_67_nl;
  wire[0:0] mem_inst_load_store_for_4_and_113_nl;
  wire[0:0] mem_inst_load_store_for_4_and_83_nl;
  wire[0:0] mem_inst_load_store_for_4_and_98_nl;
  wire[0:0] and_697_nl;
  wire[2:0] crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_8_nl;
  wire[1:0] mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_4_nl;
  wire[0:0] mem_inst_load_store_for_4_and_110_nl;
  wire[0:0] mem_inst_load_store_for_4_and_65_nl;
  wire[0:0] mem_inst_load_store_for_4_and_111_nl;
  wire[0:0] mem_inst_load_store_for_4_and_81_nl;
  wire[0:0] mem_inst_load_store_for_4_and_96_nl;
  wire[0:0] and_698_nl;
  wire[2:0] crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_6_nl;
  wire[1:0] mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_3_nl;
  wire[0:0] mem_inst_load_store_for_4_and_108_nl;
  wire[0:0] mem_inst_load_store_for_4_and_63_nl;
  wire[0:0] mem_inst_load_store_for_4_and_109_nl;
  wire[0:0] mem_inst_load_store_for_4_and_79_nl;
  wire[0:0] mem_inst_load_store_for_4_and_94_nl;
  wire[0:0] and_699_nl;
  wire[2:0] crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_4_nl;
  wire[1:0] mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_2_nl;
  wire[0:0] mem_inst_load_store_for_4_and_106_nl;
  wire[0:0] mem_inst_load_store_for_4_and_61_nl;
  wire[0:0] mem_inst_load_store_for_4_and_107_nl;
  wire[0:0] mem_inst_load_store_for_4_and_77_nl;
  wire[0:0] mem_inst_load_store_for_4_and_92_nl;
  wire[0:0] and_700_nl;
  wire[2:0] crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_2_nl;
  wire[1:0] mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_1_nl;
  wire[0:0] mem_inst_load_store_for_4_and_104_nl;
  wire[0:0] mem_inst_load_store_for_4_and_59_nl;
  wire[0:0] mem_inst_load_store_for_4_and_105_nl;
  wire[0:0] mem_inst_load_store_for_4_and_75_nl;
  wire[0:0] mem_inst_load_store_for_4_and_90_nl;
  wire[0:0] and_701_nl;
  wire[2:0] crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_nl;
  wire[1:0] mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_nl;
  wire[0:0] mem_inst_load_store_for_4_and_nl;
  wire[0:0] mem_inst_load_store_for_4_and_56_nl;
  wire[0:0] mem_inst_load_store_for_4_and_103_nl;
  wire[0:0] mem_inst_load_store_for_4_and_73_nl;
  wire[0:0] mem_inst_load_store_for_4_and_88_nl;
  wire[0:0] and_702_nl;
  wire[2:0] mem_inst_request_xbar_xbar_for_3_if_1_mux_7_nl;
  wire[2:0] mem_inst_request_xbar_xbar_for_3_if_1_mux_11_nl;
  wire[2:0] mem_inst_request_xbar_xbar_for_3_if_1_mux_15_nl;
  wire[2:0] mem_inst_request_xbar_xbar_for_3_if_1_mux_19_nl;
  wire[2:0] mem_inst_request_xbar_xbar_for_3_if_1_mux_23_nl;
  wire[2:0] mem_inst_request_xbar_xbar_for_3_if_1_mux_27_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_30_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_28_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_26_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_24_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_22_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_20_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_18_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_16_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_42_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_43_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_44_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_45_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_46_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_47_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_1_operator_3_false_operator_3_false_operator_3_false_or_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_1_operator_4_false_operator_4_false_operator_4_false_or_nl;
  wire[0:0] and_340_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_36_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_37_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_38_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_39_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_40_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_41_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_2_operator_3_false_operator_3_false_operator_3_false_or_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_2_operator_4_false_operator_4_false_operator_4_false_or_nl;
  wire[0:0] and_363_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_30_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_31_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_32_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_33_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_34_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_35_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_3_operator_3_false_operator_3_false_operator_3_false_or_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_3_operator_4_false_operator_4_false_operator_4_false_or_nl;
  wire[0:0] and_386_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_24_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_25_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_26_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_27_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_28_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_29_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_4_operator_3_false_operator_3_false_operator_3_false_or_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_4_operator_4_false_operator_4_false_operator_4_false_or_nl;
  wire[0:0] and_409_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_18_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_19_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_20_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_21_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_22_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_23_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_5_operator_3_false_operator_3_false_operator_3_false_or_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_5_operator_4_false_operator_4_false_operator_4_false_or_nl;
  wire[0:0] and_431_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_16_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_17_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_6_operator_3_false_operator_3_false_operator_3_false_or_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_6_operator_4_false_operator_4_false_operator_4_false_or_nl;
  wire[0:0] and_452_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_6_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_7_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_7_operator_3_false_operator_3_false_operator_3_false_or_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_7_operator_4_false_operator_4_false_operator_4_false_or_nl;
  wire[0:0] and_473_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_1_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_2_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_3_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_4_nl;
  wire[0:0] nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_5_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_8_operator_3_false_operator_3_false_operator_3_false_or_nl;
  wire[0:0] mem_inst_request_xbar_xbar_for_3_8_operator_4_false_operator_4_false_operator_4_false_or_nl;
  wire[0:0] and_494_nl;
  wire[0:0] while_else_while_else_or_10_nl;
  wire[0:0] while_else_while_else_or_11_nl;
  wire[0:0] while_else_while_else_or_12_nl;
  wire[0:0] while_else_while_else_or_13_nl;
  wire[0:0] while_else_while_else_or_14_nl;
  wire[0:0] while_else_while_else_or_15_nl;
  wire[0:0] while_else_while_else_or_16_nl;
  wire[0:0] while_else_while_else_or_17_nl;
  wire[2:0] mem_inst_request_xbar_xbar_for_3_if_1_mux_3_nl;
  wire[0:0] mem_inst_load_store_for_4_if_or_71_nl;
  wire[0:0] mem_inst_load_store_for_4_if_or_69_nl;
  wire[0:0] mem_inst_load_store_for_4_if_or_67_nl;
  wire[0:0] mem_inst_load_store_for_4_if_or_65_nl;
  wire[0:0] mem_inst_load_store_for_4_if_or_64_nl;
  wire[0:0] mem_inst_load_store_for_4_if_or_66_nl;
  wire[0:0] mem_inst_load_store_for_4_if_or_68_nl;
  wire[0:0] mem_inst_load_store_for_4_if_or_70_nl;
  wire[2:0] mem_inst_request_xbar_xbar_for_3_if_1_mux_31_nl;
  wire[0:0] mux_3_nl;
  wire[0:0] mux_2_nl;
  wire[0:0] mux_1_nl;
  wire[0:0] nor_45_nl;
  wire[0:0] nor_46_nl;
  wire[0:0] mux_6_nl;
  wire[0:0] mux_5_nl;
  wire[0:0] mux_4_nl;
  wire[0:0] nor_38_nl;
  wire[0:0] nor_39_nl;
  wire[0:0] nor_40_nl;
  wire[0:0] nor_41_nl;
  wire[0:0] mux_9_nl;
  wire[0:0] mux_8_nl;
  wire[0:0] mux_7_nl;
  wire[0:0] or_171_nl;
  wire[0:0] or_170_nl;
  wire[0:0] or_169_nl;
  wire[0:0] mux_12_nl;
  wire[0:0] mux_11_nl;
  wire[0:0] mux_10_nl;
  wire[0:0] nor_34_nl;
  wire[0:0] nor_35_nl;
  wire[0:0] nor_36_nl;
  wire[0:0] nor_37_nl;
  wire[0:0] mux_15_nl;
  wire[0:0] mux_14_nl;
  wire[0:0] mux_13_nl;
  wire[0:0] or_191_nl;
  wire[0:0] or_190_nl;
  wire[0:0] or_189_nl;
  wire[0:0] mux_18_nl;
  wire[0:0] mux_17_nl;
  wire[0:0] mux_16_nl;
  wire[0:0] nor_30_nl;
  wire[0:0] nor_31_nl;
  wire[0:0] nor_32_nl;
  wire[0:0] nor_33_nl;
  wire[0:0] mux_21_nl;
  wire[0:0] mux_20_nl;
  wire[0:0] mux_19_nl;
  wire[0:0] or_211_nl;
  wire[0:0] or_210_nl;
  wire[0:0] or_209_nl;
  wire[0:0] mux_24_nl;
  wire[0:0] mux_23_nl;
  wire[0:0] mux_22_nl;
  wire[0:0] nor_26_nl;
  wire[0:0] nor_27_nl;
  wire[0:0] nor_28_nl;
  wire[0:0] nor_29_nl;
  wire[0:0] mux_27_nl;
  wire[0:0] mux_26_nl;
  wire[0:0] mux_25_nl;
  wire[0:0] or_231_nl;
  wire[0:0] or_230_nl;
  wire[0:0] or_229_nl;
  wire[0:0] mux_30_nl;
  wire[0:0] mux_29_nl;
  wire[0:0] mux_28_nl;
  wire[0:0] nor_22_nl;
  wire[0:0] nor_23_nl;
  wire[0:0] nor_24_nl;
  wire[0:0] nor_25_nl;
  wire[0:0] mux_33_nl;
  wire[0:0] mux_32_nl;
  wire[0:0] mux_31_nl;
  wire[0:0] or_251_nl;
  wire[0:0] or_250_nl;
  wire[0:0] or_249_nl;
  wire[0:0] mux_36_nl;
  wire[0:0] mux_35_nl;
  wire[0:0] mux_34_nl;
  wire[0:0] nor_18_nl;
  wire[0:0] nor_19_nl;
  wire[0:0] nor_20_nl;
  wire[0:0] nor_21_nl;
  wire[0:0] mux_39_nl;
  wire[0:0] mux_38_nl;
  wire[0:0] mux_37_nl;
  wire[0:0] nor_nl;
  wire[0:0] nor_42_nl;
  wire[0:0] mux_42_nl;
  wire[0:0] mux_41_nl;
  wire[0:0] mux_40_nl;
  wire[0:0] nor_14_nl;
  wire[0:0] nor_15_nl;
  wire[0:0] nor_16_nl;
  wire[0:0] nor_17_nl;
  wire[0:0] mux_45_nl;
  wire[0:0] mux_44_nl;
  wire[0:0] mux_43_nl;
  wire[0:0] or_290_nl;
  wire[0:0] or_289_nl;
  wire[0:0] or_288_nl;
  wire[0:0] mux_48_nl;
  wire[0:0] mux_47_nl;
  wire[0:0] mux_46_nl;
  wire[0:0] nor_10_nl;
  wire[0:0] nor_11_nl;
  wire[0:0] nor_12_nl;
  wire[0:0] nor_13_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [2:0] nl_mem_inst_request_xbar_xbar_for_7_lshift_rg_s;
  assign nl_mem_inst_request_xbar_xbar_for_7_lshift_rg_s = MUX_v_3_2_2((while_req_reg_addr_sva_1[50:48]),
      3'b110, while_and_21_cse_1);
  wire [2:0] nl_mem_inst_request_xbar_xbar_for_1_lshift_rg_s;
  assign nl_mem_inst_request_xbar_xbar_for_1_lshift_rg_s = MUX_v_3_2_2((signext_3_1(~
      write_req_PopNB_mioi_return_rsc_z_mxwt)), (while_req_reg_addr_sva_1[2:0]),
      or_dcpl_40);
  wire [2:0] nl_mem_inst_request_xbar_xbar_for_8_lshift_rg_s;
  assign nl_mem_inst_request_xbar_xbar_for_8_lshift_rg_s = MUX_v_3_2_2(({{2{write_req_PopNB_mioi_return_rsc_z_mxwt}},
      write_req_PopNB_mioi_return_rsc_z_mxwt}), (while_req_reg_addr_sva_1[58:56]),
      or_dcpl_40);
  wire [2:0] nl_mem_inst_request_xbar_xbar_for_3_lshift_rg_s;
  assign nl_mem_inst_request_xbar_xbar_for_3_lshift_rg_s = MUX_v_3_2_2((while_req_reg_addr_sva_1[18:16]),
      3'b010, while_and_21_cse_1);
  wire [2:0] nl_mem_inst_request_xbar_xbar_for_5_lshift_rg_s;
  assign nl_mem_inst_request_xbar_xbar_for_5_lshift_rg_s = MUX_v_3_2_2((while_req_reg_addr_sva_1[34:32]),
      3'b100, while_and_21_cse_1);
  wire [2:0] nl_mem_inst_request_xbar_xbar_for_4_lshift_rg_s;
  assign nl_mem_inst_request_xbar_xbar_for_4_lshift_rg_s = MUX_v_3_2_2((while_req_reg_addr_sva_1[26:24]),
      3'b011, while_and_21_cse_1);
  wire [2:0] nl_mem_inst_request_xbar_xbar_for_6_lshift_rg_s;
  assign nl_mem_inst_request_xbar_xbar_for_6_lshift_rg_s = MUX_v_3_2_2((while_req_reg_addr_sva_1[42:40]),
      3'b101, while_and_21_cse_1);
  wire [2:0] nl_mem_inst_request_xbar_xbar_for_2_lshift_rg_s;
  assign nl_mem_inst_request_xbar_xbar_for_2_lshift_rg_s = MUX_v_3_2_2((while_req_reg_addr_sva_1[10:8]),
      3'b001, while_and_21_cse_1);
  wire [0:0] nl_InputSetup_MemoryRun_req_inter_PopNB_mioi_inst_req_inter_PopNB_mioi_oswt_pff;
  assign nl_InputSetup_MemoryRun_req_inter_PopNB_mioi_inst_req_inter_PopNB_mioi_oswt_pff
      = fsm_output[1];
  wire [7:0] nl_InputSetup_MemoryRun_rsp_inter_Push_mioi_inst_rsp_inter_Push_mioi_m_valids_rsc_dat_MemoryRun;
  assign nl_InputSetup_MemoryRun_rsp_inter_Push_mioi_inst_rsp_inter_Push_mioi_m_valids_rsc_dat_MemoryRun
      = {crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1_2 , crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1_dfm_1_2
      , crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1_dfm_1_2 , crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1_dfm_1_2
      , crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1_dfm_1_2 , crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1_dfm_1_2
      , crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1_dfm_1_2 , crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1_dfm_1_2};
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_6_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_5_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_4_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_3_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_2_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_1_nl;
  wire[7:0] crossbar_InputSetup_InputType_8U_8U_for_mux_nl;
  wire[7:0] mem_inst_load_store_data_out_mux_nl;
  wire [63:0] nl_InputSetup_MemoryRun_rsp_inter_Push_mioi_inst_rsp_inter_Push_mioi_m_data_rsc_dat_MemoryRun;
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_6_nl = MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
      crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
      crossbar_InputSetup_InputType_8U_8U_for_and_20_cse);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_5_nl = MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
      crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
      crossbar_InputSetup_InputType_8U_8U_for_and_20_cse);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_4_nl = MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
      crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
      crossbar_InputSetup_InputType_8U_8U_for_and_20_cse);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_3_nl = MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
      crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
      crossbar_InputSetup_InputType_8U_8U_for_and_20_cse);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_2_nl = MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
      crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
      crossbar_InputSetup_InputType_8U_8U_for_and_20_cse);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_1_nl = MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
      crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
      crossbar_InputSetup_InputType_8U_8U_for_and_20_cse);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_nl = MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
      crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
      crossbar_InputSetup_InputType_8U_8U_for_and_20_cse);
  assign mem_inst_load_store_data_out_mux_nl = MUX_v_8_2_2(mem_inst_load_store_data_out_0_lpi_1_dfm_1,
      mem_inst_load_store_data_out_0_lpi_1_dfm_2, crossbar_InputSetup_InputType_8U_8U_for_and_20_cse);
  assign nl_InputSetup_MemoryRun_rsp_inter_Push_mioi_inst_rsp_inter_Push_mioi_m_data_rsc_dat_MemoryRun
      = {(crossbar_InputSetup_InputType_8U_8U_for_mux_6_nl) , (crossbar_InputSetup_InputType_8U_8U_for_mux_5_nl)
      , (crossbar_InputSetup_InputType_8U_8U_for_mux_4_nl) , (crossbar_InputSetup_InputType_8U_8U_for_mux_3_nl)
      , (crossbar_InputSetup_InputType_8U_8U_for_mux_2_nl) , (crossbar_InputSetup_InputType_8U_8U_for_mux_1_nl)
      , (crossbar_InputSetup_InputType_8U_8U_for_mux_nl) , (mem_inst_load_store_data_out_mux_nl)};
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) mem_inst_request_xbar_xbar_for_7_lshift_rg (
      .a(while_req_reg_valids_6_lpi_1_dfm_1_mx0),
      .s(nl_mem_inst_request_xbar_xbar_for_7_lshift_rg_s[2:0]),
      .z(mem_inst_request_xbar_xbar_for_7_lshift_tmp)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) mem_inst_request_xbar_xbar_for_1_lshift_rg (
      .a(while_req_reg_valids_0_lpi_1_dfm_1_mx0),
      .s(nl_mem_inst_request_xbar_xbar_for_1_lshift_rg_s[2:0]),
      .z(mem_inst_request_xbar_xbar_for_1_lshift_tmp)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) mem_inst_request_xbar_xbar_for_8_lshift_rg (
      .a(while_req_reg_valids_7_lpi_1_dfm_1_mx0),
      .s(nl_mem_inst_request_xbar_xbar_for_8_lshift_rg_s[2:0]),
      .z(mem_inst_request_xbar_xbar_for_8_lshift_tmp)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) mem_inst_request_xbar_xbar_for_3_lshift_rg (
      .a(while_req_reg_valids_2_lpi_1_dfm_1_mx0),
      .s(nl_mem_inst_request_xbar_xbar_for_3_lshift_rg_s[2:0]),
      .z(mem_inst_request_xbar_xbar_for_3_lshift_tmp)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) mem_inst_request_xbar_xbar_for_5_lshift_rg (
      .a(while_req_reg_valids_4_lpi_1_dfm_1_mx0),
      .s(nl_mem_inst_request_xbar_xbar_for_5_lshift_rg_s[2:0]),
      .z(mem_inst_request_xbar_xbar_for_5_lshift_tmp)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) mem_inst_request_xbar_xbar_for_4_lshift_rg (
      .a(while_req_reg_valids_3_lpi_1_dfm_1_mx0),
      .s(nl_mem_inst_request_xbar_xbar_for_4_lshift_rg_s[2:0]),
      .z(mem_inst_request_xbar_xbar_for_4_lshift_tmp)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) mem_inst_request_xbar_xbar_for_6_lshift_rg (
      .a(while_req_reg_valids_5_lpi_1_dfm_1_mx0),
      .s(nl_mem_inst_request_xbar_xbar_for_6_lshift_rg_s[2:0]),
      .z(mem_inst_request_xbar_xbar_for_6_lshift_tmp)
    );
  mgc_shift_l_v5 #(.width_a(32'sd1),
  .signd_a(32'sd0),
  .width_s(32'sd3),
  .width_z(32'sd8)) mem_inst_request_xbar_xbar_for_2_lshift_rg (
      .a(while_req_reg_valids_1_lpi_1_dfm_1_mx0),
      .s(nl_mem_inst_request_xbar_xbar_for_2_lshift_rg_s[2:0]),
      .z(mem_inst_request_xbar_xbar_for_2_lshift_tmp)
    );
  InputSetup_MemoryRun_req_inter_PopNB_mioi InputSetup_MemoryRun_req_inter_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .req_inter_val(req_inter_val),
      .req_inter_rdy(req_inter_rdy),
      .req_inter_msg(req_inter_msg),
      .MemoryRun_wen(rsp_inter_Push_mioi_wen_comp),
      .req_inter_PopNB_mioi_oswt(reg_req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse),
      .MemoryRun_wten(MemoryRun_wten),
      .req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt(req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt),
      .req_inter_PopNB_mioi_data_valids_rsc_z_mxwt(req_inter_PopNB_mioi_data_valids_rsc_z_mxwt),
      .req_inter_PopNB_mioi_data_addr_rsc_z_mxwt(req_inter_PopNB_mioi_data_addr_rsc_z_mxwt),
      .req_inter_PopNB_mioi_data_data_rsc_z_mxwt(req_inter_PopNB_mioi_data_data_rsc_z_mxwt),
      .req_inter_PopNB_mioi_return_rsc_z_mxwt(req_inter_PopNB_mioi_return_rsc_z_mxwt),
      .req_inter_PopNB_mioi_oswt_pff(nl_InputSetup_MemoryRun_req_inter_PopNB_mioi_inst_req_inter_PopNB_mioi_oswt_pff[0:0]),
      .MemoryRun_wten_pff(MemoryRun_wten_iff)
    );
  InputSetup_MemoryRun_write_req_PopNB_mioi InputSetup_MemoryRun_write_req_PopNB_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .write_req_val(write_req_val),
      .write_req_rdy(write_req_rdy),
      .write_req_msg(write_req_msg),
      .MemoryRun_wen(rsp_inter_Push_mioi_wen_comp),
      .MemoryRun_wten(MemoryRun_wten),
      .write_req_PopNB_mioi_oswt(reg_write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse),
      .write_req_PopNB_mioi_data_data_data_rsc_z_mxwt(write_req_PopNB_mioi_data_data_data_rsc_z_mxwt),
      .write_req_PopNB_mioi_data_index_rsc_z_mxwt(write_req_PopNB_mioi_data_index_rsc_z_mxwt),
      .write_req_PopNB_mioi_return_rsc_z_mxwt(write_req_PopNB_mioi_return_rsc_z_mxwt),
      .write_req_PopNB_mioi_oswt_pff(and_231_rmff),
      .MemoryRun_wten_pff(MemoryRun_wten_iff)
    );
  InputSetup_MemoryRun_rsp_inter_Push_mioi InputSetup_MemoryRun_rsp_inter_Push_mioi_inst
      (
      .clk(clk),
      .rst(rst),
      .rsp_inter_val(rsp_inter_val),
      .rsp_inter_rdy(rsp_inter_rdy),
      .rsp_inter_msg(rsp_inter_msg),
      .MemoryRun_wen(rsp_inter_Push_mioi_wen_comp),
      .MemoryRun_wten(MemoryRun_wten_iff),
      .rsp_inter_Push_mioi_oswt(reg_rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse),
      .rsp_inter_Push_mioi_wen_comp(rsp_inter_Push_mioi_wen_comp),
      .rsp_inter_Push_mioi_m_valids_rsc_dat_MemoryRun(nl_InputSetup_MemoryRun_rsp_inter_Push_mioi_inst_rsp_inter_Push_mioi_m_valids_rsc_dat_MemoryRun[7:0]),
      .rsp_inter_Push_mioi_m_data_rsc_dat_MemoryRun(nl_InputSetup_MemoryRun_rsp_inter_Push_mioi_inst_rsp_inter_Push_mioi_m_data_rsc_dat_MemoryRun[63:0]),
      .rsp_inter_Push_mioi_oswt_pff(and_dcpl)
    );
  InputSetup_MemoryRun_wait_dp InputSetup_MemoryRun_wait_dp_inst (
      .clk(clk),
      .rst(rst),
      .mem_inst_banks_bank_array_impl_data0_rsc_cgo_iro(and_525_rmff),
      .mem_inst_banks_bank_array_impl_data0_rsci_data_out_d(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data0_rsci_en_d(mem_inst_banks_bank_array_impl_data0_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data1_rsc_cgo_iro(and_523_rmff),
      .mem_inst_banks_bank_array_impl_data1_rsci_data_out_d(mem_inst_banks_bank_array_impl_data1_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data1_rsci_en_d(mem_inst_banks_bank_array_impl_data1_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data2_rsc_cgo_iro(and_521_rmff),
      .mem_inst_banks_bank_array_impl_data2_rsci_data_out_d(mem_inst_banks_bank_array_impl_data2_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data2_rsci_en_d(mem_inst_banks_bank_array_impl_data2_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data3_rsc_cgo_iro(and_519_rmff),
      .mem_inst_banks_bank_array_impl_data3_rsci_data_out_d(mem_inst_banks_bank_array_impl_data3_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data3_rsci_en_d(mem_inst_banks_bank_array_impl_data3_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data4_rsc_cgo_iro(and_517_rmff),
      .mem_inst_banks_bank_array_impl_data4_rsci_data_out_d(mem_inst_banks_bank_array_impl_data4_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data4_rsci_en_d(mem_inst_banks_bank_array_impl_data4_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data5_rsc_cgo_iro(and_515_rmff),
      .mem_inst_banks_bank_array_impl_data5_rsci_data_out_d(mem_inst_banks_bank_array_impl_data5_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data5_rsci_en_d(mem_inst_banks_bank_array_impl_data5_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data6_rsc_cgo_iro(and_513_rmff),
      .mem_inst_banks_bank_array_impl_data6_rsci_data_out_d(mem_inst_banks_bank_array_impl_data6_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data6_rsci_en_d(mem_inst_banks_bank_array_impl_data6_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data7_rsc_cgo_iro(and_511_rmff),
      .mem_inst_banks_bank_array_impl_data7_rsci_data_out_d(mem_inst_banks_bank_array_impl_data7_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data7_rsci_en_d(mem_inst_banks_bank_array_impl_data7_rsci_en_d),
      .MemoryRun_wen(rsp_inter_Push_mioi_wen_comp),
      .mem_inst_banks_bank_array_impl_data0_rsc_cgo(reg_mem_inst_banks_bank_array_impl_data0_rsc_cgo_cse),
      .mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg),
      .mem_inst_banks_bank_array_impl_data1_rsc_cgo(reg_mem_inst_banks_bank_array_impl_data1_rsc_cgo_cse),
      .mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg(mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg),
      .mem_inst_banks_bank_array_impl_data2_rsc_cgo(reg_mem_inst_banks_bank_array_impl_data2_rsc_cgo_cse),
      .mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg(mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg),
      .mem_inst_banks_bank_array_impl_data3_rsc_cgo(reg_mem_inst_banks_bank_array_impl_data3_rsc_cgo_cse),
      .mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg(mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg),
      .mem_inst_banks_bank_array_impl_data4_rsc_cgo(reg_mem_inst_banks_bank_array_impl_data4_rsc_cgo_cse),
      .mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg(mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg),
      .mem_inst_banks_bank_array_impl_data5_rsc_cgo(reg_mem_inst_banks_bank_array_impl_data5_rsc_cgo_cse),
      .mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg(mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg),
      .mem_inst_banks_bank_array_impl_data6_rsc_cgo(reg_mem_inst_banks_bank_array_impl_data6_rsc_cgo_cse),
      .mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg(mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg),
      .mem_inst_banks_bank_array_impl_data7_rsc_cgo(reg_mem_inst_banks_bank_array_impl_data7_rsc_cgo_cse),
      .mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg(mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg)
    );
  InputSetup_MemoryRun_staller InputSetup_MemoryRun_staller_inst (
      .clk(clk),
      .rst(rst),
      .MemoryRun_wten(MemoryRun_wten),
      .rsp_inter_Push_mioi_wen_comp(rsp_inter_Push_mioi_wen_comp),
      .MemoryRun_wten_pff(MemoryRun_wten_iff)
    );
  InputSetup_MemoryRun_MemoryRun_fsm InputSetup_MemoryRun_MemoryRun_fsm_inst (
      .clk(clk),
      .rst(rst),
      .rsp_inter_Push_mioi_wen_comp(rsp_inter_Push_mioi_wen_comp),
      .fsm_output(fsm_output)
    );
  assign and_30_nl = and_tmp & and_685_cse & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_tmp);
  assign mem_inst_banks_read_for_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_30_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb = mem_inst_banks_read_for_mux_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_1_InputSetup_MemoryRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_30_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb = mem_inst_banks_read_for_mux_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb = mem_inst_banks_read_for_mux_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 127
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_1_InputSetup_MemoryRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_30_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb = mem_inst_banks_read_for_mux_cse;
  assign and_32_nl = and_tmp & and_685_cse & mem_inst_request_xbar_xbar_for_3_if_1_mux_tmp;
  assign mem_inst_banks_write_if_for_if_mux_cse = MUX1HOT_s_1_1_2(1'b1, and_32_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 = mem_inst_banks_write_if_for_if_mux_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_1_InputSetup_MemoryRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_32_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_1 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_1 = mem_inst_banks_write_if_for_if_mux_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 = mem_inst_banks_write_if_for_if_mux_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 147
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_1_InputSetup_MemoryRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_32_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_1 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_1 = mem_inst_banks_write_if_for_if_mux_cse;
  assign and_35_nl = and_tmp_1 & and_685_cse & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp);
  assign mem_inst_banks_read_for_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_35_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 = mem_inst_banks_read_for_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_2_InputSetup_MemoryRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_35_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_2 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_2 = mem_inst_banks_read_for_mux_4_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 = mem_inst_banks_read_for_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 127
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_2_InputSetup_MemoryRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_35_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_2 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_2 = mem_inst_banks_read_for_mux_4_cse;
  assign and_37_nl = and_tmp_1 & and_685_cse & mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp;
  assign mem_inst_banks_write_if_for_if_mux_4_cse = MUX1HOT_s_1_1_2(1'b1, and_37_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 = mem_inst_banks_write_if_for_if_mux_4_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_2_InputSetup_MemoryRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_37_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_3 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_3 = mem_inst_banks_write_if_for_if_mux_4_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 = mem_inst_banks_write_if_for_if_mux_4_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 147
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_2_InputSetup_MemoryRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_37_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_3 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_3 = mem_inst_banks_write_if_for_if_mux_4_cse;
  assign and_40_nl = and_tmp_2 & and_685_cse & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp);
  assign mem_inst_banks_read_for_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_40_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 = mem_inst_banks_read_for_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_3_InputSetup_MemoryRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_40_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_4 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_4 = mem_inst_banks_read_for_mux_8_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 = mem_inst_banks_read_for_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 127
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_3_InputSetup_MemoryRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_40_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_4 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_4 = mem_inst_banks_read_for_mux_8_cse;
  assign and_42_nl = and_tmp_2 & and_685_cse & mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp;
  assign mem_inst_banks_write_if_for_if_mux_8_cse = MUX1HOT_s_1_1_2(1'b1, and_42_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 = mem_inst_banks_write_if_for_if_mux_8_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_3_InputSetup_MemoryRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_42_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_5 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_5 = mem_inst_banks_write_if_for_if_mux_8_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 = mem_inst_banks_write_if_for_if_mux_8_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 147
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_3_InputSetup_MemoryRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_42_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_5 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_5 = mem_inst_banks_write_if_for_if_mux_8_cse;
  assign and_45_nl = and_tmp_3 & and_685_cse & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp);
  assign mem_inst_banks_read_for_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_45_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 = mem_inst_banks_read_for_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_4_InputSetup_MemoryRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_45_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_6 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_6 = mem_inst_banks_read_for_mux_12_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 = mem_inst_banks_read_for_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 127
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_4_InputSetup_MemoryRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_45_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_6 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_6 = mem_inst_banks_read_for_mux_12_cse;
  assign and_47_nl = and_tmp_3 & and_685_cse & mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp;
  assign mem_inst_banks_write_if_for_if_mux_12_cse = MUX1HOT_s_1_1_2(1'b1, and_47_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 = mem_inst_banks_write_if_for_if_mux_12_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_4_InputSetup_MemoryRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_47_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_7 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_7 = mem_inst_banks_write_if_for_if_mux_12_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 = mem_inst_banks_write_if_for_if_mux_12_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 147
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_4_InputSetup_MemoryRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_47_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_7 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_7 = mem_inst_banks_write_if_for_if_mux_12_cse;
  assign and_50_nl = and_tmp_4 & and_685_cse & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp);
  assign mem_inst_banks_read_for_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_50_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 = mem_inst_banks_read_for_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_5_InputSetup_MemoryRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_50_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_8 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_8 = mem_inst_banks_read_for_mux_16_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 = mem_inst_banks_read_for_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 127
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_5_InputSetup_MemoryRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_50_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_8 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_8 = mem_inst_banks_read_for_mux_16_cse;
  assign and_52_nl = and_tmp_4 & and_685_cse & mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp;
  assign mem_inst_banks_write_if_for_if_mux_16_cse = MUX1HOT_s_1_1_2(1'b1, and_52_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 = mem_inst_banks_write_if_for_if_mux_16_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_5_InputSetup_MemoryRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_52_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_9 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_9 = mem_inst_banks_write_if_for_if_mux_16_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 = mem_inst_banks_write_if_for_if_mux_16_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 147
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_5_InputSetup_MemoryRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_52_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_9 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_9 = mem_inst_banks_write_if_for_if_mux_16_cse;
  assign and_55_nl = and_tmp_5 & and_685_cse & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp);
  assign mem_inst_banks_read_for_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_55_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 = mem_inst_banks_read_for_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_6_InputSetup_MemoryRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_55_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_10 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_10 = mem_inst_banks_read_for_mux_20_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 = mem_inst_banks_read_for_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 127
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_6_InputSetup_MemoryRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_55_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_10 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_10 = mem_inst_banks_read_for_mux_20_cse;
  assign and_57_nl = and_tmp_5 & and_685_cse & mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp;
  assign mem_inst_banks_write_if_for_if_mux_20_cse = MUX1HOT_s_1_1_2(1'b1, and_57_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 = mem_inst_banks_write_if_for_if_mux_20_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_6_InputSetup_MemoryRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_57_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_11 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_11 = mem_inst_banks_write_if_for_if_mux_20_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 = mem_inst_banks_write_if_for_if_mux_20_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 147
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_6_InputSetup_MemoryRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_57_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_11 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_11 = mem_inst_banks_write_if_for_if_mux_20_cse;
  assign and_60_nl = and_tmp_6 & and_685_cse & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp);
  assign mem_inst_banks_read_for_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_60_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 = mem_inst_banks_read_for_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_7_InputSetup_MemoryRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_60_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_12 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_12 = mem_inst_banks_read_for_mux_24_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 = mem_inst_banks_read_for_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 127
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_7_InputSetup_MemoryRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_60_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_12 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_12 = mem_inst_banks_read_for_mux_24_cse;
  assign and_62_nl = and_tmp_6 & and_685_cse & mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp;
  assign mem_inst_banks_write_if_for_if_mux_24_cse = MUX1HOT_s_1_1_2(1'b1, and_62_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 = mem_inst_banks_write_if_for_if_mux_24_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_7_InputSetup_MemoryRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_62_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_13 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_13 = mem_inst_banks_write_if_for_if_mux_24_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 = mem_inst_banks_write_if_for_if_mux_24_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 147
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_7_InputSetup_MemoryRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_62_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_13 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_13 = mem_inst_banks_write_if_for_if_mux_24_cse;
  assign and_65_nl = and_tmp_7 & and_685_cse & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_28_tmp);
  assign mem_inst_banks_read_for_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_65_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 = mem_inst_banks_read_for_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 126
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_8_InputSetup_MemoryRun_mem_array_h_ln126_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_65_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_14 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_14 = mem_inst_banks_read_for_mux_28_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 = mem_inst_banks_read_for_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 127
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_8_InputSetup_MemoryRun_mem_array_h_ln127_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_65_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_14 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_14 = mem_inst_banks_read_for_mux_28_cse;
  assign and_67_nl = and_tmp_7 & and_685_cse & mem_inst_request_xbar_xbar_for_3_if_1_mux_28_tmp;
  assign mem_inst_banks_write_if_for_if_mux_28_cse = MUX1HOT_s_1_1_2(1'b1, and_67_nl);
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 = mem_inst_banks_write_if_for_if_mux_28_cse;
  // assert(bank_sel<NumBanks && "bank_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 146
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_8_InputSetup_MemoryRun_mem_array_h_ln146_assert_bank_sel_lt_NumBanks_and_bank_index_out_of_bounds : assert always ( rst && and_67_nl -> pbank_sel_NumBanks_bank_index_out_of_bounds_prb_15 );
  assign pbank_sel_NumBanks_bank_index_out_of_bounds_ctrl_prb_15 = mem_inst_banks_write_if_for_if_mux_28_cse;
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 = mem_inst_banks_write_if_for_if_mux_28_cse;
  // assert(idx<NumEntriesPerBank && "local_index_out_of_bounds") - ../../../matchlib/cmod/include/mem_array.h: line 147
  // psl default clock = (posedge clk);
  // psl mem_inst_banks_load_store_for_8_InputSetup_MemoryRun_mem_array_h_ln147_assert_idx_lt_NumEntriesPerBank_and_local_index_out_of_bounds : assert always ( rst && and_67_nl -> pidx_NumEntriesPerBank_local_index_out_of_bounds_prb_15 );
  assign pidx_NumEntriesPerBank_local_index_out_of_bounds_ctrl_prb_15 = mem_inst_banks_write_if_for_if_mux_28_cse;
  assign and_511_rmff = ((and_tmp_7 & and_685_cse) | (and_dcpl_1 & mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1))
      & (fsm_output[1]);
  assign and_513_rmff = ((and_tmp_6 & and_685_cse) | (and_dcpl_1 & mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1))
      & (fsm_output[1]);
  assign and_515_rmff = ((and_tmp_5 & and_685_cse) | (and_dcpl_1 & mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1))
      & (fsm_output[1]);
  assign and_517_rmff = ((and_tmp_4 & and_685_cse) | (and_dcpl_1 & mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1))
      & (fsm_output[1]);
  assign and_519_rmff = ((and_tmp_3 & and_685_cse) | (and_dcpl_1 & mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1))
      & (fsm_output[1]);
  assign and_521_rmff = ((and_tmp_2 & and_685_cse) | (and_dcpl_1 & mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1))
      & (fsm_output[1]);
  assign and_523_rmff = ((and_tmp_1 & and_685_cse) | (and_dcpl_1 & mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1))
      & (fsm_output[1]);
  assign and_525_rmff = ((and_tmp & and_685_cse) | (and_dcpl_1 & mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1))
      & (fsm_output[1]);
  assign and_231_rmff = reg_req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse
      & (~ req_inter_PopNB_mioi_return_rsc_z_mxwt);
  assign crossbar_InputSetup_InputType_8U_8U_for_aelse_and_8_cse = rsp_inter_Push_mioi_wen_comp
      & or_dcpl_1 & and_dcpl_1;
  assign or_2_nl = while_lor_lpi_1_dfm_st_1 | (~ nor_tmp_1);
  assign mux_nl = MUX_s_1_2_2(and_dcpl_1, (or_2_nl), and_685_cse);
  assign crossbar_InputSetup_InputType_8U_8U_for_and_7_cse = rsp_inter_Push_mioi_wen_comp
      & (~ (fsm_output[0])) & (~ (mux_nl));
  assign crossbar_InputSetup_InputType_8U_8U_for_aelse_and_16_cse = rsp_inter_Push_mioi_wen_comp
      & nor_tmp_1;
  assign while_and_itm = rsp_inter_Push_mioi_wen_comp & while_stage_0_4;
  assign mem_inst_request_xbar_xbar_for_3_and_cse = rsp_inter_Push_mioi_wen_comp
      & and_685_cse;
  assign while_oelse_and_1_cse = rsp_inter_Push_mioi_wen_comp & while_stage_0_3;
  assign while_req_reg_addr_and_cse = rsp_inter_Push_mioi_wen_comp & reg_req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse;
  assign mem_inst_request_xbar_arbiters_next_and_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~((mem_inst_request_xbar_xbar_for_2_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[0])
      | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[0])
      | (~ and_dcpl_122))) | or_dcpl_12));
  assign mem_inst_request_xbar_arbiters_next_and_7_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~((~ and_dcpl_131) | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[1])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[1])
      | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[1])
      | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[1]))) | or_dcpl_12));
  assign mem_inst_request_xbar_arbiters_next_and_14_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~((mem_inst_request_xbar_xbar_for_5_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[2])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[2])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[2])
      | (~ and_dcpl_134))) | or_dcpl_12));
  assign mem_inst_request_xbar_arbiters_next_and_21_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~((mem_inst_request_xbar_xbar_for_5_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[3])
      | (~ and_dcpl_144) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[3])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[3])))
      | or_dcpl_12));
  assign mem_inst_request_xbar_arbiters_next_and_28_cse = rsp_inter_Push_mioi_wen_comp
      & (~(((~ (mem_inst_request_xbar_xbar_for_4_lshift_tmp[4])) & (~ (mem_inst_request_xbar_xbar_for_5_lshift_tmp[4]))
      & and_dcpl_151 & (~ (mem_inst_request_xbar_xbar_for_2_lshift_tmp[4])) & (~
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[4])) & and_dcpl_148) | or_dcpl_12));
  assign mem_inst_request_xbar_arbiters_next_and_35_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~((mem_inst_request_xbar_xbar_for_2_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[5])
      | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[5])
      | (~ and_dcpl_157))) | or_dcpl_12));
  assign mem_inst_request_xbar_arbiters_next_and_42_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~((~ and_dcpl_167) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[6])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[6])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[6]))) | or_dcpl_12));
  assign operator_15_false_and_cse = rsp_inter_Push_mioi_wen_comp & (~((~((mem_inst_request_xbar_xbar_for_3_lshift_tmp[7])
      | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[7])
      | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[7]) | (~ and_dcpl_171))) | or_dcpl_12));
  assign crossbar_InputSetup_InputType_8U_8U_for_aelse_and_cse = rsp_inter_Push_mioi_wen_comp
      & (~ or_dcpl_12);
  assign mem_inst_load_store_for_4_if_and_104_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~ and_tmp_1) | or_dcpl_12 | mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp));
  assign mem_inst_load_store_for_4_if_and_108_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~ and_tmp_2) | or_dcpl_12 | mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp));
  assign mem_inst_load_store_for_4_if_and_112_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~ and_tmp_3) | or_dcpl_12 | mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp));
  assign mem_inst_load_store_for_4_if_and_116_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~ and_tmp_4) | or_dcpl_12 | mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp));
  assign mem_inst_load_store_for_4_if_and_120_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~ and_tmp_5) | or_dcpl_12 | mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp));
  assign mem_inst_load_store_for_4_if_and_124_cse = rsp_inter_Push_mioi_wen_comp
      & (~((~ and_tmp_6) | or_dcpl_12 | mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp));
  assign mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1
      = mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | (mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_15) | (mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_15) | (mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_15) | (mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_15) | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  assign mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1
      = mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | (mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_14) | (mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_14) | (mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_14) | (mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_14) | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  assign mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1
      = mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | (mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_13) | (mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_13) | (mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_13) | (mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_13) | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  assign mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1
      = mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | (mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_12) | (mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_12) | (mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_12) | (mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_12) | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  assign mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1
      = mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | (mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_11) | (mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_11) | (mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_11) | (mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_11) | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  assign mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1
      = mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | (mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_10) | (mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_10) | (mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_10) | (mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_10) | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  assign mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1
      = mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | (mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_9) | (mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_9) | (mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_9) | (mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_9) | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  assign mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1
      = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | (mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_8) | (mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_8) | (mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_8) | (mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_8) | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7;
  assign while_if_1_while_if_1_or_tmp = write_req_PopNB_mioi_return_rsc_z_mxwt |
      while_asn_mdf_sva_1;
  assign and_687_tmp = (~(mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1 & mem_inst_load_store_for_4_if_and_tmp_8_sva_1))
      & mem_inst_load_store_valid_src_7_lpi_1_dfm_7_mx0;
  assign crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_14_nl
      = MUX_v_3_2_2(3'b000, ({{2{mem_inst_load_store_valid_src_7_lpi_1_dfm_7_mx0}},
      mem_inst_load_store_valid_src_7_lpi_1_dfm_7_mx0}), mem_inst_load_store_for_4_if_and_tmp_8_sva_1);
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_7_nl
      = MUX_v_2_2_2((signext_2_1(~ mem_inst_load_store_for_4_if_and_tmp_sva_2)),
      2'b01, mem_inst_load_store_for_4_and_55_cse_1);
  assign mem_inst_load_store_for_4_and_116_nl = (~(mem_inst_load_store_for_4_and_7_tmp_1
      | mem_inst_load_store_for_4_and_15_tmp_1)) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_23_m1c_1
      & and_687_tmp;
  assign mem_inst_load_store_for_4_and_71_nl = mem_inst_load_store_for_4_and_7_tmp_1
      & (~ mem_inst_load_store_for_4_and_15_tmp_1) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_23_m1c_1
      & and_687_tmp;
  assign mem_inst_load_store_for_4_and_117_nl = mem_inst_load_store_for_4_and_15_tmp_1
      & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_23_m1c_1 & and_687_tmp;
  assign mem_inst_load_store_for_4_and_87_nl = mem_inst_load_store_for_4_and_23_tmp_1
      & (~ mem_inst_load_store_for_4_and_31_tmp_1) & (~ mem_inst_load_store_for_4_and_39_tmp_1)
      & and_687_tmp;
  assign mem_inst_load_store_for_4_and_102_nl = mem_inst_load_store_for_4_and_31_tmp_1
      & (~ mem_inst_load_store_for_4_and_39_tmp_1) & and_687_tmp;
  assign and_695_nl = mem_inst_load_store_for_4_and_39_tmp_1 & and_687_tmp;
  assign crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_1 = MUX1HOT_v_3_7_2((crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_14_nl),
      (signext_3_2(mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_7_nl)),
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, {(~ and_687_tmp) , (mem_inst_load_store_for_4_and_116_nl)
      , (mem_inst_load_store_for_4_and_71_nl) , (mem_inst_load_store_for_4_and_117_nl)
      , (mem_inst_load_store_for_4_and_87_nl) , (mem_inst_load_store_for_4_and_102_nl)
      , (and_695_nl)});
  assign and_688_tmp = (~(mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1 & mem_inst_load_store_for_4_if_and_tmp_9_sva_1))
      & mem_inst_load_store_valid_src_6_lpi_1_dfm_7_mx0;
  assign crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_12_nl
      = MUX_v_3_2_2(3'b000, ({{2{mem_inst_load_store_valid_src_6_lpi_1_dfm_7_mx0}},
      mem_inst_load_store_valid_src_6_lpi_1_dfm_7_mx0}), mem_inst_load_store_for_4_if_and_tmp_9_sva_1);
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_6_nl
      = MUX_v_2_2_2((signext_2_1(~ mem_inst_load_store_for_4_if_and_tmp_1_sva_2)),
      2'b01, mem_inst_load_store_for_4_and_53_cse_1);
  assign mem_inst_load_store_for_4_and_114_nl = (~(mem_inst_load_store_for_4_and_6_tmp_1
      | mem_inst_load_store_for_4_and_14_tmp_1)) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_22_m1c_1
      & and_688_tmp;
  assign mem_inst_load_store_for_4_and_69_nl = mem_inst_load_store_for_4_and_6_tmp_1
      & (~ mem_inst_load_store_for_4_and_14_tmp_1) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_22_m1c_1
      & and_688_tmp;
  assign mem_inst_load_store_for_4_and_115_nl = mem_inst_load_store_for_4_and_14_tmp_1
      & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_22_m1c_1 & and_688_tmp;
  assign mem_inst_load_store_for_4_and_85_nl = mem_inst_load_store_for_4_and_22_tmp_1
      & (~ mem_inst_load_store_for_4_and_30_tmp_1) & (~ mem_inst_load_store_for_4_and_38_tmp_1)
      & and_688_tmp;
  assign mem_inst_load_store_for_4_and_100_nl = mem_inst_load_store_for_4_and_30_tmp_1
      & (~ mem_inst_load_store_for_4_and_38_tmp_1) & and_688_tmp;
  assign and_696_nl = mem_inst_load_store_for_4_and_38_tmp_1 & and_688_tmp;
  assign crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_1 = MUX1HOT_v_3_7_2((crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_12_nl),
      (signext_3_2(mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_6_nl)),
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, {(~ and_688_tmp) , (mem_inst_load_store_for_4_and_114_nl)
      , (mem_inst_load_store_for_4_and_69_nl) , (mem_inst_load_store_for_4_and_115_nl)
      , (mem_inst_load_store_for_4_and_85_nl) , (mem_inst_load_store_for_4_and_100_nl)
      , (and_696_nl)});
  assign and_689_tmp = (~(mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1 & mem_inst_load_store_for_4_if_and_tmp_10_sva_1))
      & mem_inst_load_store_valid_src_5_lpi_1_dfm_7_mx0;
  assign crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_10_nl
      = MUX_v_3_2_2(3'b000, ({{2{mem_inst_load_store_valid_src_5_lpi_1_dfm_7_mx0}},
      mem_inst_load_store_valid_src_5_lpi_1_dfm_7_mx0}), mem_inst_load_store_for_4_if_and_tmp_10_sva_1);
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_5_nl
      = MUX_v_2_2_2((signext_2_1(~ mem_inst_load_store_for_4_if_and_tmp_2_sva_2)),
      2'b01, mem_inst_load_store_for_4_and_51_cse_1);
  assign mem_inst_load_store_for_4_and_112_nl = (~(mem_inst_load_store_for_4_and_5_tmp_1
      | mem_inst_load_store_for_4_and_13_tmp_1)) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_21_m1c_1
      & and_689_tmp;
  assign mem_inst_load_store_for_4_and_67_nl = mem_inst_load_store_for_4_and_5_tmp_1
      & (~ mem_inst_load_store_for_4_and_13_tmp_1) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_21_m1c_1
      & and_689_tmp;
  assign mem_inst_load_store_for_4_and_113_nl = mem_inst_load_store_for_4_and_13_tmp_1
      & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_21_m1c_1 & and_689_tmp;
  assign mem_inst_load_store_for_4_and_83_nl = mem_inst_load_store_for_4_and_21_tmp_1
      & (~ mem_inst_load_store_for_4_and_29_tmp_1) & (~ mem_inst_load_store_for_4_and_37_tmp_1)
      & and_689_tmp;
  assign mem_inst_load_store_for_4_and_98_nl = mem_inst_load_store_for_4_and_29_tmp_1
      & (~ mem_inst_load_store_for_4_and_37_tmp_1) & and_689_tmp;
  assign and_697_nl = mem_inst_load_store_for_4_and_37_tmp_1 & and_689_tmp;
  assign crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_1 = MUX1HOT_v_3_7_2((crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_10_nl),
      (signext_3_2(mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_5_nl)),
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, {(~ and_689_tmp) , (mem_inst_load_store_for_4_and_112_nl)
      , (mem_inst_load_store_for_4_and_67_nl) , (mem_inst_load_store_for_4_and_113_nl)
      , (mem_inst_load_store_for_4_and_83_nl) , (mem_inst_load_store_for_4_and_98_nl)
      , (and_697_nl)});
  assign and_690_tmp = (~(mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1 & mem_inst_load_store_for_4_if_and_tmp_11_sva_1))
      & mem_inst_load_store_valid_src_4_lpi_1_dfm_7_mx0;
  assign crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_8_nl
      = MUX_v_3_2_2(3'b000, ({{2{mem_inst_load_store_valid_src_4_lpi_1_dfm_7_mx0}},
      mem_inst_load_store_valid_src_4_lpi_1_dfm_7_mx0}), mem_inst_load_store_for_4_if_and_tmp_11_sva_1);
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_4_nl
      = MUX_v_2_2_2((signext_2_1(~ mem_inst_load_store_for_4_if_and_tmp_3_sva_2)),
      2'b01, mem_inst_load_store_for_4_and_49_cse_1);
  assign mem_inst_load_store_for_4_and_110_nl = (~(mem_inst_load_store_for_4_and_4_tmp_1
      | mem_inst_load_store_for_4_and_12_tmp_1)) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_20_m1c_1
      & and_690_tmp;
  assign mem_inst_load_store_for_4_and_65_nl = mem_inst_load_store_for_4_and_4_tmp_1
      & (~ mem_inst_load_store_for_4_and_12_tmp_1) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_20_m1c_1
      & and_690_tmp;
  assign mem_inst_load_store_for_4_and_111_nl = mem_inst_load_store_for_4_and_12_tmp_1
      & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_20_m1c_1 & and_690_tmp;
  assign mem_inst_load_store_for_4_and_81_nl = mem_inst_load_store_for_4_and_20_tmp_1
      & (~ mem_inst_load_store_for_4_and_28_tmp_1) & (~ mem_inst_load_store_for_4_and_36_tmp_1)
      & and_690_tmp;
  assign mem_inst_load_store_for_4_and_96_nl = mem_inst_load_store_for_4_and_28_tmp_1
      & (~ mem_inst_load_store_for_4_and_36_tmp_1) & and_690_tmp;
  assign and_698_nl = mem_inst_load_store_for_4_and_36_tmp_1 & and_690_tmp;
  assign crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_1 = MUX1HOT_v_3_7_2((crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_8_nl),
      (signext_3_2(mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_4_nl)),
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, {(~ and_690_tmp) , (mem_inst_load_store_for_4_and_110_nl)
      , (mem_inst_load_store_for_4_and_65_nl) , (mem_inst_load_store_for_4_and_111_nl)
      , (mem_inst_load_store_for_4_and_81_nl) , (mem_inst_load_store_for_4_and_96_nl)
      , (and_698_nl)});
  assign and_691_tmp = (~(mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1 & mem_inst_load_store_for_4_if_and_tmp_12_sva_1))
      & mem_inst_load_store_valid_src_3_lpi_1_dfm_7_mx0;
  assign crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_6_nl
      = MUX_v_3_2_2(3'b000, ({{2{mem_inst_load_store_valid_src_3_lpi_1_dfm_7_mx0}},
      mem_inst_load_store_valid_src_3_lpi_1_dfm_7_mx0}), mem_inst_load_store_for_4_if_and_tmp_12_sva_1);
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_3_nl
      = MUX_v_2_2_2((signext_2_1(~ mem_inst_load_store_for_4_if_and_tmp_4_sva_2)),
      2'b01, mem_inst_load_store_for_4_and_47_cse_1);
  assign mem_inst_load_store_for_4_and_108_nl = (~(mem_inst_load_store_for_4_and_3_tmp_1
      | mem_inst_load_store_for_4_and_11_tmp_1)) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_19_m1c_1
      & and_691_tmp;
  assign mem_inst_load_store_for_4_and_63_nl = mem_inst_load_store_for_4_and_3_tmp_1
      & (~ mem_inst_load_store_for_4_and_11_tmp_1) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_19_m1c_1
      & and_691_tmp;
  assign mem_inst_load_store_for_4_and_109_nl = mem_inst_load_store_for_4_and_11_tmp_1
      & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_19_m1c_1 & and_691_tmp;
  assign mem_inst_load_store_for_4_and_79_nl = mem_inst_load_store_for_4_and_19_tmp_1
      & (~ mem_inst_load_store_for_4_and_27_tmp_1) & (~ mem_inst_load_store_for_4_and_35_tmp_1)
      & and_691_tmp;
  assign mem_inst_load_store_for_4_and_94_nl = mem_inst_load_store_for_4_and_27_tmp_1
      & (~ mem_inst_load_store_for_4_and_35_tmp_1) & and_691_tmp;
  assign and_699_nl = mem_inst_load_store_for_4_and_35_tmp_1 & and_691_tmp;
  assign crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_1 = MUX1HOT_v_3_7_2((crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_6_nl),
      (signext_3_2(mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_3_nl)),
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, {(~ and_691_tmp) , (mem_inst_load_store_for_4_and_108_nl)
      , (mem_inst_load_store_for_4_and_63_nl) , (mem_inst_load_store_for_4_and_109_nl)
      , (mem_inst_load_store_for_4_and_79_nl) , (mem_inst_load_store_for_4_and_94_nl)
      , (and_699_nl)});
  assign and_692_tmp = (~(mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1 & mem_inst_load_store_for_4_if_and_tmp_13_sva_1))
      & mem_inst_load_store_valid_src_2_lpi_1_dfm_7_mx0;
  assign crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_4_nl
      = MUX_v_3_2_2(3'b000, ({{2{mem_inst_load_store_valid_src_2_lpi_1_dfm_7_mx0}},
      mem_inst_load_store_valid_src_2_lpi_1_dfm_7_mx0}), mem_inst_load_store_for_4_if_and_tmp_13_sva_1);
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_2_nl
      = MUX_v_2_2_2((signext_2_1(~ mem_inst_load_store_for_4_if_and_tmp_5_sva_2)),
      2'b01, mem_inst_load_store_for_4_and_45_cse_1);
  assign mem_inst_load_store_for_4_and_106_nl = (~(mem_inst_load_store_for_4_and_2_tmp_1
      | mem_inst_load_store_for_4_and_10_tmp_1)) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_18_m1c_1
      & and_692_tmp;
  assign mem_inst_load_store_for_4_and_61_nl = mem_inst_load_store_for_4_and_2_tmp_1
      & (~ mem_inst_load_store_for_4_and_10_tmp_1) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_18_m1c_1
      & and_692_tmp;
  assign mem_inst_load_store_for_4_and_107_nl = mem_inst_load_store_for_4_and_10_tmp_1
      & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_18_m1c_1 & and_692_tmp;
  assign mem_inst_load_store_for_4_and_77_nl = mem_inst_load_store_for_4_and_18_tmp_1
      & (~ mem_inst_load_store_for_4_and_26_tmp_1) & (~ mem_inst_load_store_for_4_and_34_tmp_1)
      & and_692_tmp;
  assign mem_inst_load_store_for_4_and_92_nl = mem_inst_load_store_for_4_and_26_tmp_1
      & (~ mem_inst_load_store_for_4_and_34_tmp_1) & and_692_tmp;
  assign and_700_nl = mem_inst_load_store_for_4_and_34_tmp_1 & and_692_tmp;
  assign crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_1 = MUX1HOT_v_3_7_2((crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_4_nl),
      (signext_3_2(mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_2_nl)),
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, {(~ and_692_tmp) , (mem_inst_load_store_for_4_and_106_nl)
      , (mem_inst_load_store_for_4_and_61_nl) , (mem_inst_load_store_for_4_and_107_nl)
      , (mem_inst_load_store_for_4_and_77_nl) , (mem_inst_load_store_for_4_and_92_nl)
      , (and_700_nl)});
  assign and_693_tmp = (~(mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1 & mem_inst_load_store_for_4_if_and_tmp_14_sva_1))
      & mem_inst_load_store_valid_src_1_lpi_1_dfm_7_mx0;
  assign crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_2_nl
      = MUX_v_3_2_2(3'b000, ({{2{mem_inst_load_store_valid_src_1_lpi_1_dfm_7_mx0}},
      mem_inst_load_store_valid_src_1_lpi_1_dfm_7_mx0}), mem_inst_load_store_for_4_if_and_tmp_14_sva_1);
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_1_nl
      = MUX_v_2_2_2((signext_2_1(~ mem_inst_load_store_for_4_if_and_tmp_6_sva_2)),
      2'b01, mem_inst_load_store_for_4_and_43_cse_1);
  assign mem_inst_load_store_for_4_and_104_nl = (~(mem_inst_load_store_for_4_and_1_tmp_1
      | mem_inst_load_store_for_4_and_9_tmp_1)) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_17_m1c_1
      & and_693_tmp;
  assign mem_inst_load_store_for_4_and_59_nl = mem_inst_load_store_for_4_and_1_tmp_1
      & (~ mem_inst_load_store_for_4_and_9_tmp_1) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_17_m1c_1
      & and_693_tmp;
  assign mem_inst_load_store_for_4_and_105_nl = mem_inst_load_store_for_4_and_9_tmp_1
      & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_17_m1c_1 & and_693_tmp;
  assign mem_inst_load_store_for_4_and_75_nl = mem_inst_load_store_for_4_and_17_tmp_1
      & (~ mem_inst_load_store_for_4_and_25_tmp_1) & (~ mem_inst_load_store_for_4_and_33_tmp_1)
      & and_693_tmp;
  assign mem_inst_load_store_for_4_and_90_nl = mem_inst_load_store_for_4_and_25_tmp_1
      & (~ mem_inst_load_store_for_4_and_33_tmp_1) & and_693_tmp;
  assign and_701_nl = mem_inst_load_store_for_4_and_33_tmp_1 & and_693_tmp;
  assign crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_1 = MUX1HOT_v_3_7_2((crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_2_nl),
      (signext_3_2(mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_1_nl)),
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, {(~ and_693_tmp) , (mem_inst_load_store_for_4_and_104_nl)
      , (mem_inst_load_store_for_4_and_59_nl) , (mem_inst_load_store_for_4_and_105_nl)
      , (mem_inst_load_store_for_4_and_75_nl) , (mem_inst_load_store_for_4_and_90_nl)
      , (and_701_nl)});
  assign and_694_tmp = (or_dcpl_137 | (~ mem_inst_load_store_for_4_if_and_tmp_15_sva_1))
      & mem_inst_load_store_valid_src_0_lpi_1_dfm_7_mx0;
  assign crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_nl
      = MUX_v_3_2_2(3'b000, ({{2{mem_inst_load_store_valid_src_0_lpi_1_dfm_7_mx0}},
      mem_inst_load_store_valid_src_0_lpi_1_dfm_7_mx0}), mem_inst_load_store_for_4_if_and_tmp_15_sva_1);
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_nl
      = MUX_v_2_2_2((signext_2_1(~ mem_inst_load_store_for_4_if_and_tmp_7_sva_2)),
      2'b01, mem_inst_load_store_for_4_and_41_cse_1);
  assign mem_inst_load_store_for_4_and_nl = (~(mem_inst_load_store_for_4_and_tmp_1
      | mem_inst_load_store_for_4_and_8_tmp_1)) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_16_m1c_1
      & and_694_tmp;
  assign mem_inst_load_store_for_4_and_56_nl = mem_inst_load_store_for_4_and_tmp_1
      & (~ mem_inst_load_store_for_4_and_8_tmp_1) & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_16_m1c_1
      & and_694_tmp;
  assign mem_inst_load_store_for_4_and_103_nl = mem_inst_load_store_for_4_and_8_tmp_1
      & mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_16_m1c_1 & and_694_tmp;
  assign mem_inst_load_store_for_4_and_73_nl = mem_inst_load_store_for_4_and_16_tmp_1
      & (~ mem_inst_load_store_for_4_and_24_tmp_1) & (~ mem_inst_load_store_for_4_and_32_tmp_1)
      & and_694_tmp;
  assign mem_inst_load_store_for_4_and_88_nl = mem_inst_load_store_for_4_and_24_tmp_1
      & (~ mem_inst_load_store_for_4_and_32_tmp_1) & and_694_tmp;
  assign and_702_nl = mem_inst_load_store_for_4_and_32_tmp_1 & and_694_tmp;
  assign crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_1 = MUX1HOT_v_3_7_2((crossbar_InputSetup_InputType_8U_8U_for_crossbar_InputSetup_InputType_8U_8U_for_and_nl),
      (signext_3_2(mem_inst_load_store_for_4_mem_inst_load_store_for_4_mem_inst_load_store_for_4_mux_nl)),
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, {(~ and_694_tmp) , (mem_inst_load_store_for_4_and_nl)
      , (mem_inst_load_store_for_4_and_56_nl) , (mem_inst_load_store_for_4_and_103_nl)
      , (mem_inst_load_store_for_4_and_73_nl) , (mem_inst_load_store_for_4_and_88_nl)
      , (and_702_nl)});
  assign mem_inst_load_store_for_4_if_and_stg_1_0_1_sva_mx0w0 = ~((mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx0w0[1:0]!=2'b00));
  assign mem_inst_load_store_for_4_if_and_stg_1_0_1_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_0_1_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_0_1_sva, or_dcpl_24);
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_7_nl = MUX_v_3_8_2(3'b000, 3'b001,
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_2_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_2_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_2_sva_1});
  assign mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx0w0 =
      MUX_v_3_2_2(3'b000, (mem_inst_request_xbar_xbar_for_3_if_1_mux_7_nl), mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1);
  assign mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2 =
      MUX_s_1_2_2((mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx0w0[2]),
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_ftd, or_dcpl_24);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_1_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx0w0[1:0]==2'b01);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_1_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_1_1_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_1_1_sva, or_dcpl_24);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_1_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx0w0[1:0]==2'b10);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_1_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_2_1_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_2_1_sva, or_dcpl_24);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_1_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx0w0[1:0]==2'b11);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_1_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_3_1_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_3_1_sva, or_dcpl_24);
  assign mem_inst_load_store_for_4_if_and_stg_1_0_2_sva_mx0w0 = ~((mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx0w0[1:0]!=2'b00));
  assign mem_inst_load_store_for_4_if_and_stg_1_0_2_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_0_2_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_0_2_sva, or_dcpl_27);
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_11_nl = MUX_v_3_8_2(3'b000, 3'b001,
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_3_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_3_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_3_sva_1});
  assign mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx0w0 =
      MUX_v_3_2_2(3'b000, (mem_inst_request_xbar_xbar_for_3_if_1_mux_11_nl), mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1);
  assign mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2 =
      MUX_s_1_2_2((mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx0w0[2]),
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_ftd, or_dcpl_27);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_2_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx0w0[1:0]==2'b01);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_2_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_1_2_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_1_2_sva, or_dcpl_27);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_2_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx0w0[1:0]==2'b10);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_2_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_2_2_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_2_2_sva, or_dcpl_27);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_2_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx0w0[1:0]==2'b11);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_2_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_3_2_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_3_2_sva, or_dcpl_27);
  assign mem_inst_load_store_for_4_if_and_stg_1_0_3_sva_mx0w0 = ~((mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx0w0[1:0]!=2'b00));
  assign mem_inst_load_store_for_4_if_and_stg_1_0_3_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_0_3_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_0_3_sva, or_dcpl_30);
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_15_nl = MUX_v_3_8_2(3'b000, 3'b001,
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_4_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_4_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_4_sva_1});
  assign mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx0w0 =
      MUX_v_3_2_2(3'b000, (mem_inst_request_xbar_xbar_for_3_if_1_mux_15_nl), mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1);
  assign mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2 =
      MUX_s_1_2_2((mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx0w0[2]),
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_ftd, or_dcpl_30);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_3_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx0w0[1:0]==2'b01);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_3_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_1_3_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_1_3_sva, or_dcpl_30);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_3_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx0w0[1:0]==2'b10);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_3_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_2_3_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_2_3_sva, or_dcpl_30);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_3_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx0w0[1:0]==2'b11);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_3_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_3_3_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_3_3_sva, or_dcpl_30);
  assign mem_inst_load_store_for_4_if_and_stg_1_0_4_sva_mx0w0 = ~((mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx0w0[1:0]!=2'b00));
  assign mem_inst_load_store_for_4_if_and_stg_1_0_4_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_0_4_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_0_4_sva, or_dcpl_33);
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_19_nl = MUX_v_3_8_2(3'b000, 3'b001,
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_5_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_5_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_5_sva_1});
  assign mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx0w0 =
      MUX_v_3_2_2(3'b000, (mem_inst_request_xbar_xbar_for_3_if_1_mux_19_nl), mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1);
  assign mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2 =
      MUX_s_1_2_2((mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx0w0[2]),
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_ftd, or_dcpl_33);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_4_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx0w0[1:0]==2'b01);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_4_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_1_4_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_1_4_sva, or_dcpl_33);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_4_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx0w0[1:0]==2'b10);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_4_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_2_4_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_2_4_sva, or_dcpl_33);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_4_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx0w0[1:0]==2'b11);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_4_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_3_4_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_3_4_sva, or_dcpl_33);
  assign mem_inst_load_store_for_4_if_and_stg_1_0_5_sva_mx0w0 = ~((mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx0w0[1:0]!=2'b00));
  assign mem_inst_load_store_for_4_if_and_stg_1_0_5_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_0_5_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_0_5_sva, or_dcpl_36);
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_23_nl = MUX_v_3_8_2(3'b000, 3'b001,
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_6_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_6_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_6_sva_1});
  assign mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx0w0 =
      MUX_v_3_2_2(3'b000, (mem_inst_request_xbar_xbar_for_3_if_1_mux_23_nl), mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1);
  assign mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2 =
      MUX_s_1_2_2((mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx0w0[2]),
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_ftd, or_dcpl_36);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_5_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx0w0[1:0]==2'b01);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_5_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_1_5_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_1_5_sva, or_dcpl_36);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_5_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx0w0[1:0]==2'b10);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_5_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_2_5_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_2_5_sva, or_dcpl_36);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_5_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx0w0[1:0]==2'b11);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_5_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_3_5_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_3_5_sva, or_dcpl_36);
  assign mem_inst_load_store_for_4_if_and_stg_1_0_6_sva_mx0w0 = ~((mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx0w0[1:0]!=2'b00));
  assign mem_inst_load_store_for_4_if_and_stg_1_0_6_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_0_6_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_0_6_sva, or_dcpl_39);
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_27_nl = MUX_v_3_8_2(3'b000, 3'b001,
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_7_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_7_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_7_sva_1});
  assign mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx0w0 =
      MUX_v_3_2_2(3'b000, (mem_inst_request_xbar_xbar_for_3_if_1_mux_27_nl), mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1);
  assign mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2 =
      MUX_s_1_2_2((mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx0w0[2]),
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_ftd, or_dcpl_39);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_6_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx0w0[1:0]==2'b01);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_6_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_1_6_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_1_6_sva, or_dcpl_39);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_6_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx0w0[1:0]==2'b10);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_6_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_2_6_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_2_6_sva, or_dcpl_39);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_6_sva_mx0w0 = (mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx0w0[1:0]==2'b11);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_6_sva_mx1 = MUX_s_1_2_2(mem_inst_load_store_for_4_if_and_stg_1_3_6_sva_mx0w0,
      mem_inst_load_store_for_4_if_and_stg_1_3_6_sva, or_dcpl_39);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_30_nl = MUX_v_8_8_2(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg, crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2
      = MUX_v_8_2_2(8'b00000000, (crossbar_InputSetup_InputType_8U_8U_for_mux_30_nl),
      crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_28_nl = MUX_v_8_8_2(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg, crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2
      = MUX_v_8_2_2(8'b00000000, (crossbar_InputSetup_InputType_8U_8U_for_mux_28_nl),
      crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_26_nl = MUX_v_8_8_2(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg, crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2
      = MUX_v_8_2_2(8'b00000000, (crossbar_InputSetup_InputType_8U_8U_for_mux_26_nl),
      crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_24_nl = MUX_v_8_8_2(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg, crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2
      = MUX_v_8_2_2(8'b00000000, (crossbar_InputSetup_InputType_8U_8U_for_mux_24_nl),
      crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_22_nl = MUX_v_8_8_2(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg, crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2
      = MUX_v_8_2_2(8'b00000000, (crossbar_InputSetup_InputType_8U_8U_for_mux_22_nl),
      crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_20_nl = MUX_v_8_8_2(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg, crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2
      = MUX_v_8_2_2(8'b00000000, (crossbar_InputSetup_InputType_8U_8U_for_mux_20_nl),
      crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_18_nl = MUX_v_8_8_2(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg, crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2
      = MUX_v_8_2_2(8'b00000000, (crossbar_InputSetup_InputType_8U_8U_for_mux_18_nl),
      crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1_dfm_2);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_16_nl = MUX_v_8_8_2(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data1_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data2_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data3_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data4_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data5_rsci_data_out_d_oreg, mem_inst_banks_bank_array_impl_data6_rsci_data_out_d_oreg,
      mem_inst_banks_bank_array_impl_data7_rsci_data_out_d_oreg, crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_2);
  assign mem_inst_load_store_data_out_0_lpi_1_dfm_2 = MUX_v_8_2_2(8'b00000000, (crossbar_InputSetup_InputType_8U_8U_for_mux_16_nl),
      crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1_dfm_2);
  assign while_req_reg_data_0_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((write_req_PopNB_mioi_data_data_data_rsc_z_mxwt[7:0]),
      (while_req_reg_data_sva_1[7:0]), or_dcpl_40);
  assign while_req_reg_data_1_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((write_req_PopNB_mioi_data_data_data_rsc_z_mxwt[15:8]),
      (while_req_reg_data_sva_1[15:8]), or_dcpl_40);
  assign while_req_reg_data_2_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((write_req_PopNB_mioi_data_data_data_rsc_z_mxwt[23:16]),
      (while_req_reg_data_sva_1[23:16]), or_dcpl_40);
  assign while_req_reg_data_3_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((write_req_PopNB_mioi_data_data_data_rsc_z_mxwt[31:24]),
      (while_req_reg_data_sva_1[31:24]), or_dcpl_40);
  assign while_req_reg_data_4_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((write_req_PopNB_mioi_data_data_data_rsc_z_mxwt[39:32]),
      (while_req_reg_data_sva_1[39:32]), or_dcpl_40);
  assign while_req_reg_data_5_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((write_req_PopNB_mioi_data_data_data_rsc_z_mxwt[47:40]),
      (while_req_reg_data_sva_1[47:40]), or_dcpl_40);
  assign while_req_reg_data_6_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((write_req_PopNB_mioi_data_data_data_rsc_z_mxwt[55:48]),
      (while_req_reg_data_sva_1[55:48]), or_dcpl_40);
  assign while_req_reg_data_7_lpi_1_dfm_1_mx0 = MUX_v_8_2_2((write_req_PopNB_mioi_data_data_data_rsc_z_mxwt[63:56]),
      (while_req_reg_data_sva_1[63:56]), or_dcpl_40);
  assign while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0 = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      (while_req_reg_addr_sva_1[7:3]), or_dcpl_40);
  assign while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0 = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      (while_req_reg_addr_sva_1[15:11]), or_dcpl_40);
  assign while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0 = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      (while_req_reg_addr_sva_1[23:19]), or_dcpl_40);
  assign while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0 = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      (while_req_reg_addr_sva_1[31:27]), or_dcpl_40);
  assign while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0 = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      (while_req_reg_addr_sva_1[39:35]), or_dcpl_40);
  assign while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0 = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      (while_req_reg_addr_sva_1[47:43]), or_dcpl_40);
  assign while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0 = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      (while_req_reg_addr_sva_1[55:51]), or_dcpl_40);
  assign while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0 = MUX_v_5_2_2(write_req_PopNB_mioi_data_index_rsc_z_mxwt,
      (while_req_reg_addr_sva_1[63:59]), or_dcpl_40);
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_tmp = MUX_s_1_8_2(mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_lpi_1_dfm_1, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_1_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_1_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_1_sva_1});
  assign one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_1_sva_1 =
      mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_1_sva_1 =
      mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_1_sva_1 =
      mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1 = while_req_reg_type_val_lpi_1_dfm_2
      & while_req_reg_valids_0_lpi_1_dfm_1_mx0;
  assign mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1 = while_req_reg_type_val_lpi_1_dfm_2
      & while_req_reg_valids_1_lpi_1_dfm_1_mx0;
  assign mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1 = while_req_reg_type_val_lpi_1_dfm_2
      & while_req_reg_valids_2_lpi_1_dfm_1_mx0;
  assign mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1 = while_req_reg_type_val_lpi_1_dfm_2
      & while_req_reg_valids_3_lpi_1_dfm_1_mx0;
  assign mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1 = while_req_reg_type_val_lpi_1_dfm_2
      & while_req_reg_valids_4_lpi_1_dfm_1_mx0;
  assign mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1 = while_req_reg_type_val_lpi_1_dfm_2
      & while_req_reg_valids_5_lpi_1_dfm_1_mx0;
  assign mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1 = while_req_reg_type_val_lpi_1_dfm_2
      & while_req_reg_valids_6_lpi_1_dfm_1_mx0;
  assign mem_inst_compute_bank_request_for_land_lpi_1_dfm_1 = while_req_reg_type_val_lpi_1_dfm_2
      & while_req_reg_valids_7_lpi_1_dfm_1_mx0;
  assign Arbiter_8U_Roundrobin_pick_unequal_tmp_8 = (mem_inst_request_xbar_xbar_for_8_lshift_tmp[0])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[0])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[0])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[0])
      | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[0]);
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0 & operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl
      = Arbiter_8U_Roundrobin_pick_priority_13_1_sva_1 & (~ Arbiter_8U_Roundrobin_pick_priority_14_1_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_42_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1) & and_dcpl_185;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_43_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1 & and_dcpl_185;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_44_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1)
      & and_dcpl_189;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_45_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1 &
      and_dcpl_189;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_46_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1)
      & and_dcpl_190;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_47_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1 &
      and_dcpl_190;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2((nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl),
      Arbiter_8U_Roundrobin_pick_priority_9_1_sva_1, Arbiter_8U_Roundrobin_pick_priority_11_1_sva_1,
      (mem_inst_request_xbar_xbar_for_7_lshift_tmp[0]), (mem_inst_request_xbar_xbar_for_1_lshift_tmp[0]),
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[0]), (mem_inst_request_xbar_xbar_for_5_lshift_tmp[0]),
      {or_dcpl_42 , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_42_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_43_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_44_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_45_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_46_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_47_nl)});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_priority_14_1_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1,
      {or_dcpl_42 , and_dcpl_185 , and_dcpl_189 , and_dcpl_190});
  assign mem_inst_request_xbar_xbar_for_3_1_operator_3_false_operator_3_false_operator_3_false_or_nl
      = Arbiter_8U_Roundrobin_pick_priority_14_1_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_1_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_12_1_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_1_operator_4_false_operator_4_false_operator_4_false_or_nl
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[0])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[0]);
  assign and_340_nl = or_dcpl_52 & or_dcpl_51 & or_dcpl_50 & or_dcpl_49 & or_dcpl_45
      & or_dcpl_44 & or_dcpl_43;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0
      = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_3_1_operator_3_false_operator_3_false_operator_3_false_or_nl),
      (mem_inst_request_xbar_xbar_for_3_1_operator_4_false_operator_4_false_operator_4_false_or_nl),
      and_340_nl);
  assign Arbiter_8U_Roundrobin_pick_priority_9_1_sva_1 = mem_inst_request_xbar_arbiters_next_0_2_sva
      & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_priority_11_1_sva_1 = mem_inst_request_xbar_arbiters_next_0_4_sva
      & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[0]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_1_sva_1 = Arbiter_8U_Roundrobin_pick_priority_11_1_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_1_sva_1;
  assign Arbiter_8U_Roundrobin_pick_priority_10_1_sva_1 = mem_inst_request_xbar_arbiters_next_0_3_sva
      & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_priority_13_1_sva_1 = mem_inst_request_xbar_arbiters_next_0_6_sva
      & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_priority_14_1_sva_1 = mem_inst_request_xbar_arbiters_next_0_7_sva
      & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[0]);
  assign Arbiter_8U_Roundrobin_pick_priority_12_1_sva_1 = mem_inst_request_xbar_arbiters_next_0_5_sva
      & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[0]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_1_sva_1
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[0]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_1_sva_1
      = (mem_inst_request_xbar_xbar_for_5_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[0]);
  assign mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      = mem_inst_request_xbar_arbiters_next_0_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[0]);
  assign operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1 = Arbiter_8U_Roundrobin_pick_priority_14_1_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_13_1_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_1_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_1_sva_1 | Arbiter_8U_Roundrobin_pick_priority_10_1_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_1_sva_1 | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp = MUX_s_1_8_2(mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_lpi_1_dfm_1, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_2_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_2_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_2_sva_1});
  assign one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_2_sva_1 =
      mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_2_sva_1 =
      mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_2_sva_1 =
      mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign Arbiter_8U_Roundrobin_pick_unequal_tmp_9 = (mem_inst_request_xbar_xbar_for_8_lshift_tmp[1])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[1])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[1])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[1])
      | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[1]);
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      = mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      = mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      = mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      = mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      = mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      = mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_1 & operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_1 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl
      = Arbiter_8U_Roundrobin_pick_priority_13_2_sva_1 & (~ Arbiter_8U_Roundrobin_pick_priority_14_2_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_36_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1) & and_dcpl_206;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_37_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1 & and_dcpl_206;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_38_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1)
      & and_dcpl_210;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_39_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1 &
      and_dcpl_210;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_40_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1)
      & and_dcpl_213;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_41_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1 &
      and_dcpl_213;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2((nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl),
      Arbiter_8U_Roundrobin_pick_priority_9_2_sva_1, Arbiter_8U_Roundrobin_pick_priority_11_2_sva_1,
      (mem_inst_request_xbar_xbar_for_7_lshift_tmp[1]), (mem_inst_request_xbar_xbar_for_1_lshift_tmp[1]),
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[1]), (mem_inst_request_xbar_xbar_for_5_lshift_tmp[1]),
      {or_dcpl_54 , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_36_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_37_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_38_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_39_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_40_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_41_nl)});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_2_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_priority_14_2_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1,
      {or_dcpl_54 , and_dcpl_206 , and_dcpl_210 , and_dcpl_213});
  assign mem_inst_request_xbar_xbar_for_3_2_operator_3_false_operator_3_false_operator_3_false_or_nl
      = Arbiter_8U_Roundrobin_pick_priority_14_2_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_2_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_12_2_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_2_operator_4_false_operator_4_false_operator_4_false_or_nl
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[1])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[1]);
  assign and_363_nl = or_dcpl_57 & or_dcpl_56 & or_dcpl_64 & or_dcpl_63 & or_dcpl_62
      & or_dcpl_61 & or_dcpl_55;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_3_2_operator_3_false_operator_3_false_operator_3_false_or_nl),
      (mem_inst_request_xbar_xbar_for_3_2_operator_4_false_operator_4_false_operator_4_false_or_nl),
      and_363_nl);
  assign Arbiter_8U_Roundrobin_pick_priority_9_2_sva_1 = mem_inst_request_xbar_arbiters_next_1_2_sva
      & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_priority_11_2_sva_1 = mem_inst_request_xbar_arbiters_next_1_4_sva
      & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[1]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_priority_11_2_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_2_sva_1;
  assign Arbiter_8U_Roundrobin_pick_priority_10_2_sva_1 = mem_inst_request_xbar_arbiters_next_1_3_sva
      & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_priority_13_2_sva_1 = mem_inst_request_xbar_arbiters_next_1_6_sva
      & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_priority_14_2_sva_1 = mem_inst_request_xbar_arbiters_next_1_7_sva
      & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[1]);
  assign Arbiter_8U_Roundrobin_pick_priority_12_2_sva_1 = mem_inst_request_xbar_arbiters_next_1_5_sva
      & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[1]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_2_sva_1
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[1]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_2_sva_1
      = (mem_inst_request_xbar_xbar_for_5_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[1]);
  assign mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      = mem_inst_request_xbar_arbiters_next_1_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[1]);
  assign operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1 = Arbiter_8U_Roundrobin_pick_priority_14_2_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_13_2_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_2_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_2_sva_1 | Arbiter_8U_Roundrobin_pick_priority_10_2_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_2_sva_1 | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp = MUX_s_1_8_2(mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_lpi_1_dfm_1, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_3_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_3_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_3_sva_1});
  assign one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_3_sva_1 =
      mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_3_sva_1 =
      mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_3_sva_1 =
      mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign Arbiter_8U_Roundrobin_pick_unequal_tmp_10 = (mem_inst_request_xbar_xbar_for_8_lshift_tmp[2])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[2])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[2])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[2])
      | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[2]);
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      = mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      = mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      = mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      = mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      = mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      = mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_2 & operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_2 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl
      = Arbiter_8U_Roundrobin_pick_priority_13_3_sva_1 & (~ Arbiter_8U_Roundrobin_pick_priority_14_3_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_30_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1) & and_dcpl_229;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_31_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1 & and_dcpl_229;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_32_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1)
      & and_dcpl_233;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_33_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1 &
      and_dcpl_233;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_34_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1)
      & and_dcpl_236;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_35_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1 &
      and_dcpl_236;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2((nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl),
      Arbiter_8U_Roundrobin_pick_priority_9_3_sva_1, Arbiter_8U_Roundrobin_pick_priority_11_3_sva_1,
      (mem_inst_request_xbar_xbar_for_7_lshift_tmp[2]), (mem_inst_request_xbar_xbar_for_1_lshift_tmp[2]),
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[2]), (mem_inst_request_xbar_xbar_for_5_lshift_tmp[2]),
      {or_dcpl_66 , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_30_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_31_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_32_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_33_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_34_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_35_nl)});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_3_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_priority_14_3_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1,
      {or_dcpl_66 , and_dcpl_229 , and_dcpl_233 , and_dcpl_236});
  assign mem_inst_request_xbar_xbar_for_3_3_operator_3_false_operator_3_false_operator_3_false_or_nl
      = Arbiter_8U_Roundrobin_pick_priority_14_3_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_3_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_12_3_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_3_operator_4_false_operator_4_false_operator_4_false_or_nl
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[2])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[2]);
  assign and_386_nl = or_dcpl_76 & or_dcpl_75 & or_dcpl_74 & or_dcpl_69 & or_dcpl_68
      & or_dcpl_73 & or_dcpl_67;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0
      = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_3_3_operator_3_false_operator_3_false_operator_3_false_or_nl),
      (mem_inst_request_xbar_xbar_for_3_3_operator_4_false_operator_4_false_operator_4_false_or_nl),
      and_386_nl);
  assign Arbiter_8U_Roundrobin_pick_priority_9_3_sva_1 = mem_inst_request_xbar_arbiters_next_2_2_sva
      & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_priority_11_3_sva_1 = mem_inst_request_xbar_arbiters_next_2_4_sva
      & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[2]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_priority_11_3_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_3_sva_1;
  assign Arbiter_8U_Roundrobin_pick_priority_10_3_sva_1 = mem_inst_request_xbar_arbiters_next_2_3_sva
      & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_priority_13_3_sva_1 = mem_inst_request_xbar_arbiters_next_2_6_sva
      & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_priority_14_3_sva_1 = mem_inst_request_xbar_arbiters_next_2_7_sva
      & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[2]);
  assign Arbiter_8U_Roundrobin_pick_priority_12_3_sva_1 = mem_inst_request_xbar_arbiters_next_2_5_sva
      & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[2]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_3_sva_1
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[2]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_3_sva_1
      = (mem_inst_request_xbar_xbar_for_5_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[2]);
  assign mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      = mem_inst_request_xbar_arbiters_next_2_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[2]);
  assign operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1 = Arbiter_8U_Roundrobin_pick_priority_14_3_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_13_3_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_3_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_3_sva_1 | Arbiter_8U_Roundrobin_pick_priority_10_3_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_3_sva_1 | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp = MUX_s_1_8_2(mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_lpi_1_dfm_1, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_4_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_4_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_4_sva_1});
  assign one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_4_sva_1 =
      mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_4_sva_1 =
      mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_4_sva_1 =
      mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign Arbiter_8U_Roundrobin_pick_unequal_tmp_11 = (mem_inst_request_xbar_xbar_for_8_lshift_tmp[3])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[3])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[3])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[3])
      | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[3]);
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_3 & operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_3 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_3 & operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_3 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_3 & operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_3 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_3 & operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_3 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_3 & operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_3 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_3 & operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_3 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_3 & operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_3 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl
      = Arbiter_8U_Roundrobin_pick_priority_13_4_sva_1 & (~ Arbiter_8U_Roundrobin_pick_priority_14_4_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_24_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1) & and_dcpl_252;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_25_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1 & and_dcpl_252;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_26_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1)
      & and_dcpl_256;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_27_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1 &
      and_dcpl_256;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_28_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1)
      & and_dcpl_259;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_29_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1 &
      and_dcpl_259;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2((nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl),
      Arbiter_8U_Roundrobin_pick_priority_9_4_sva_1, Arbiter_8U_Roundrobin_pick_priority_11_4_sva_1,
      (mem_inst_request_xbar_xbar_for_7_lshift_tmp[3]), (mem_inst_request_xbar_xbar_for_1_lshift_tmp[3]),
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[3]), (mem_inst_request_xbar_xbar_for_5_lshift_tmp[3]),
      {or_dcpl_78 , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_24_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_25_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_26_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_27_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_28_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_29_nl)});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_4_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_priority_14_4_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1,
      {or_dcpl_78 , and_dcpl_252 , and_dcpl_256 , and_dcpl_259});
  assign mem_inst_request_xbar_xbar_for_3_4_operator_3_false_operator_3_false_operator_3_false_or_nl
      = Arbiter_8U_Roundrobin_pick_priority_14_4_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_4_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_12_4_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_4_operator_4_false_operator_4_false_operator_4_false_or_nl
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[3])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[3]);
  assign and_409_nl = or_dcpl_88 & or_dcpl_87 & or_dcpl_81 & or_dcpl_80 & or_dcpl_86
      & or_dcpl_79 & or_dcpl_85;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0
      = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_3_4_operator_3_false_operator_3_false_operator_3_false_or_nl),
      (mem_inst_request_xbar_xbar_for_3_4_operator_4_false_operator_4_false_operator_4_false_or_nl),
      and_409_nl);
  assign Arbiter_8U_Roundrobin_pick_priority_9_4_sva_1 = mem_inst_request_xbar_arbiters_next_3_2_sva
      & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_priority_11_4_sva_1 = mem_inst_request_xbar_arbiters_next_3_4_sva
      & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[3]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_priority_11_4_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_4_sva_1;
  assign Arbiter_8U_Roundrobin_pick_priority_10_4_sva_1 = mem_inst_request_xbar_arbiters_next_3_3_sva
      & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_priority_13_4_sva_1 = mem_inst_request_xbar_arbiters_next_3_6_sva
      & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_priority_14_4_sva_1 = mem_inst_request_xbar_arbiters_next_3_7_sva
      & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[3]);
  assign Arbiter_8U_Roundrobin_pick_priority_12_4_sva_1 = mem_inst_request_xbar_arbiters_next_3_5_sva
      & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[3]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_4_sva_1
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[3]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_4_sva_1
      = (mem_inst_request_xbar_xbar_for_5_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[3]);
  assign mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      = mem_inst_request_xbar_arbiters_next_3_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[3]);
  assign operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1 = Arbiter_8U_Roundrobin_pick_priority_14_4_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_13_4_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_4_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_4_sva_1 | Arbiter_8U_Roundrobin_pick_priority_10_4_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_4_sva_1 | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp = MUX_s_1_8_2(mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_lpi_1_dfm_1, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_5_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_5_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_5_sva_1});
  assign one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_5_sva_1 =
      mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_5_sva_1 =
      mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_5_sva_1 =
      mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign Arbiter_8U_Roundrobin_pick_unequal_tmp_12 = (mem_inst_request_xbar_xbar_for_8_lshift_tmp[4])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[4])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[4])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[4])
      | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[4]);
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_4 & operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_4 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_4 & operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_4 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_4 & operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_4 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_4 & operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_4 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_4 & operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_4 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_4 & operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_4 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_4 & operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_4 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl
      = Arbiter_8U_Roundrobin_pick_priority_13_5_sva_1 & (~ Arbiter_8U_Roundrobin_pick_priority_14_5_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_18_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1) & and_dcpl_275;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_19_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1 & and_dcpl_275;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_20_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1)
      & and_dcpl_279;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_21_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1 &
      and_dcpl_279;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_22_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1)
      & and_dcpl_281;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_23_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1 &
      and_dcpl_281;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2((nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl),
      Arbiter_8U_Roundrobin_pick_priority_9_5_sva_1, Arbiter_8U_Roundrobin_pick_priority_11_5_sva_1,
      (mem_inst_request_xbar_xbar_for_7_lshift_tmp[4]), (mem_inst_request_xbar_xbar_for_1_lshift_tmp[4]),
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[4]), (mem_inst_request_xbar_xbar_for_5_lshift_tmp[4]),
      {or_dcpl_90 , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_18_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_19_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_20_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_21_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_22_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_23_nl)});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_5_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_priority_14_5_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1,
      {or_dcpl_90 , and_dcpl_275 , and_dcpl_279 , and_dcpl_281});
  assign mem_inst_request_xbar_xbar_for_3_5_operator_3_false_operator_3_false_operator_3_false_or_nl
      = Arbiter_8U_Roundrobin_pick_priority_14_5_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_5_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_12_5_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_5_operator_4_false_operator_4_false_operator_4_false_or_nl
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[4])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[4]);
  assign and_431_nl = or_dcpl_100 & or_dcpl_99 & or_dcpl_93 & or_dcpl_92 & or_dcpl_98
      & or_dcpl_97 & or_dcpl_91;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0
      = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_3_5_operator_3_false_operator_3_false_operator_3_false_or_nl),
      (mem_inst_request_xbar_xbar_for_3_5_operator_4_false_operator_4_false_operator_4_false_or_nl),
      and_431_nl);
  assign Arbiter_8U_Roundrobin_pick_priority_9_5_sva_1 = mem_inst_request_xbar_arbiters_next_4_2_sva
      & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_priority_11_5_sva_1 = mem_inst_request_xbar_arbiters_next_4_4_sva
      & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[4]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_priority_11_5_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_5_sva_1;
  assign Arbiter_8U_Roundrobin_pick_priority_10_5_sva_1 = mem_inst_request_xbar_arbiters_next_4_3_sva
      & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_priority_13_5_sva_1 = mem_inst_request_xbar_arbiters_next_4_6_sva
      & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_priority_14_5_sva_1 = mem_inst_request_xbar_arbiters_next_4_7_sva
      & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[4]);
  assign Arbiter_8U_Roundrobin_pick_priority_12_5_sva_1 = mem_inst_request_xbar_arbiters_next_4_5_sva
      & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[4]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_5_sva_1
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[4]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_5_sva_1
      = (mem_inst_request_xbar_xbar_for_5_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[4]);
  assign mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      = mem_inst_request_xbar_arbiters_next_4_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[4]);
  assign operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1 = Arbiter_8U_Roundrobin_pick_priority_14_5_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_13_5_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_5_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_5_sva_1 | Arbiter_8U_Roundrobin_pick_priority_10_5_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_5_sva_1 | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp = MUX_s_1_8_2(mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_lpi_1_dfm_1, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_6_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_6_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_6_sva_1});
  assign one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_6_sva_1 =
      mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_6_sva_1 =
      mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_6_sva_1 =
      mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign Arbiter_8U_Roundrobin_pick_unequal_tmp_13 = (mem_inst_request_xbar_xbar_for_8_lshift_tmp[5])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[5])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[5])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[5])
      | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[5]);
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_5 & operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_5 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_5 & operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_5 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_5 & operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_5 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_5 & operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_5 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_5 & operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_5 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_5 & operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_5 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_5 & operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_5 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl
      = Arbiter_8U_Roundrobin_pick_priority_13_6_sva_1 & (~ Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1) & and_dcpl_297;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1 & and_dcpl_297;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1)
      & and_dcpl_301;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1 &
      and_dcpl_301;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_16_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1)
      & and_dcpl_302;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_17_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1 &
      and_dcpl_302;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2((nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl),
      Arbiter_8U_Roundrobin_pick_priority_9_6_sva_1, Arbiter_8U_Roundrobin_pick_priority_11_6_sva_1,
      (mem_inst_request_xbar_xbar_for_7_lshift_tmp[5]), (mem_inst_request_xbar_xbar_for_1_lshift_tmp[5]),
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[5]), (mem_inst_request_xbar_xbar_for_5_lshift_tmp[5]),
      {or_dcpl_102 , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_12_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_13_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_16_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_17_nl)});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_6_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1,
      {or_dcpl_102 , and_dcpl_297 , and_dcpl_301 , and_dcpl_302});
  assign mem_inst_request_xbar_xbar_for_3_6_operator_3_false_operator_3_false_operator_3_false_or_nl
      = Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_6_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_12_6_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_6_operator_4_false_operator_4_false_operator_4_false_or_nl
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[5])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[5]);
  assign and_452_nl = or_dcpl_112 & or_dcpl_111 & or_dcpl_110 & or_dcpl_109 & or_dcpl_105
      & or_dcpl_104 & or_dcpl_103;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0
      = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_3_6_operator_3_false_operator_3_false_operator_3_false_or_nl),
      (mem_inst_request_xbar_xbar_for_3_6_operator_4_false_operator_4_false_operator_4_false_or_nl),
      and_452_nl);
  assign Arbiter_8U_Roundrobin_pick_priority_9_6_sva_1 = mem_inst_request_xbar_arbiters_next_5_2_sva
      & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_priority_11_6_sva_1 = mem_inst_request_xbar_arbiters_next_5_4_sva
      & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[5]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_priority_11_6_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_6_sva_1;
  assign Arbiter_8U_Roundrobin_pick_priority_10_6_sva_1 = mem_inst_request_xbar_arbiters_next_5_3_sva
      & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_priority_13_6_sva_1 = mem_inst_request_xbar_arbiters_next_5_6_sva
      & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1 = mem_inst_request_xbar_arbiters_next_5_7_sva
      & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[5]);
  assign Arbiter_8U_Roundrobin_pick_priority_12_6_sva_1 = mem_inst_request_xbar_arbiters_next_5_5_sva
      & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[5]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_6_sva_1
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[5]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_6_sva_1
      = (mem_inst_request_xbar_xbar_for_5_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[5]);
  assign mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      = mem_inst_request_xbar_arbiters_next_5_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[5]);
  assign operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1 = Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_13_6_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_6_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_6_sva_1 | Arbiter_8U_Roundrobin_pick_priority_10_6_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_6_sva_1 | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp = MUX_s_1_8_2(mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_lpi_1_dfm_1, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_7_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_7_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_7_sva_1});
  assign one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_7_sva_1 =
      mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_7_sva_1 =
      mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_7_sva_1 =
      mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign Arbiter_8U_Roundrobin_pick_unequal_tmp_14 = (mem_inst_request_xbar_xbar_for_8_lshift_tmp[6])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[6])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[6])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[6])
      | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[6]);
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_6 & operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_6 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_6 & operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_6 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_6 & operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_6 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_6 & operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_6 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_6 & operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_6 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_6 & operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_6 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_6 & operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_6 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl
      = Arbiter_8U_Roundrobin_pick_priority_13_7_sva_1 & (~ Arbiter_8U_Roundrobin_pick_priority_14_7_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_6_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1) & and_dcpl_318;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_7_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1 & and_dcpl_318;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1)
      & and_dcpl_322;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1 &
      and_dcpl_322;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1)
      & and_dcpl_323;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1 &
      and_dcpl_323;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2((nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_14_nl),
      Arbiter_8U_Roundrobin_pick_priority_9_7_sva_1, Arbiter_8U_Roundrobin_pick_priority_11_7_sva_1,
      (mem_inst_request_xbar_xbar_for_7_lshift_tmp[6]), (mem_inst_request_xbar_xbar_for_1_lshift_tmp[6]),
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[6]), (mem_inst_request_xbar_xbar_for_5_lshift_tmp[6]),
      {or_dcpl_114 , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_6_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_7_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_8_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_9_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_10_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_11_nl)});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_7_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_priority_14_7_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1,
      {or_dcpl_114 , and_dcpl_318 , and_dcpl_322 , and_dcpl_323});
  assign mem_inst_request_xbar_xbar_for_3_7_operator_3_false_operator_3_false_operator_3_false_or_nl
      = Arbiter_8U_Roundrobin_pick_priority_14_7_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_7_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_12_7_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_7_operator_4_false_operator_4_false_operator_4_false_or_nl
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[6])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[6]);
  assign and_473_nl = or_dcpl_117 & or_dcpl_116 & or_dcpl_115 & or_dcpl_124 & or_dcpl_123
      & or_dcpl_122 & or_dcpl_121;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0
      = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_3_7_operator_3_false_operator_3_false_operator_3_false_or_nl),
      (mem_inst_request_xbar_xbar_for_3_7_operator_4_false_operator_4_false_operator_4_false_or_nl),
      and_473_nl);
  assign Arbiter_8U_Roundrobin_pick_priority_9_7_sva_1 = mem_inst_request_xbar_arbiters_next_6_2_sva
      & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_priority_11_7_sva_1 = mem_inst_request_xbar_arbiters_next_6_4_sva
      & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[6]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_priority_11_7_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_7_sva_1;
  assign Arbiter_8U_Roundrobin_pick_priority_10_7_sva_1 = mem_inst_request_xbar_arbiters_next_6_3_sva
      & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_priority_13_7_sva_1 = mem_inst_request_xbar_arbiters_next_6_6_sva
      & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_priority_14_7_sva_1 = mem_inst_request_xbar_arbiters_next_6_7_sva
      & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[6]);
  assign Arbiter_8U_Roundrobin_pick_priority_12_7_sva_1 = mem_inst_request_xbar_arbiters_next_6_5_sva
      & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[6]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_7_sva_1
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[6]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_7_sva_1
      = (mem_inst_request_xbar_xbar_for_5_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[6]);
  assign mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1
      = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      = mem_inst_request_xbar_arbiters_next_6_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[6]);
  assign operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1 = Arbiter_8U_Roundrobin_pick_priority_14_7_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_13_7_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_7_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_7_sva_1 | Arbiter_8U_Roundrobin_pick_priority_10_7_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_7_sva_1 | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_28_tmp = MUX_s_1_8_2(mem_inst_compute_bank_request_for_land_1_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_2_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_3_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_4_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_5_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_6_lpi_1_dfm_1, mem_inst_compute_bank_request_for_land_7_lpi_1_dfm_1,
      mem_inst_compute_bank_request_for_land_lpi_1_dfm_1, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_sva_1});
  assign one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_sva_1 = mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_sva_1 = mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_sva_1 = mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6;
  assign Arbiter_8U_Roundrobin_pick_unequal_tmp_15 = (mem_inst_request_xbar_xbar_for_8_lshift_tmp[7])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[7])
      | (mem_inst_request_xbar_xbar_for_5_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[7])
      | (mem_inst_request_xbar_xbar_for_3_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_2_lshift_tmp[7])
      | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[7]);
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_7 & operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_7 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_7 & operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_7 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_7 & operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_7 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_7 & operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_7 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_7 & operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_7 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_7 & operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_7 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1));
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      = (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_7 & operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1)
      | (Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_7 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1));
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl
      = Arbiter_8U_Roundrobin_pick_priority_13_sva_1 & (~ Arbiter_8U_Roundrobin_pick_priority_14_sva_1);
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_nl
      = (~ operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1) & and_dcpl_339;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_1_nl
      = operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1 & and_dcpl_339;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_2_nl
      = (~ operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1)
      & and_dcpl_343;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_3_nl
      = operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1 & and_dcpl_343;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_4_nl
      = (~ operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1)
      & and_dcpl_344;
  assign nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_5_nl
      = operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1 & and_dcpl_344;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_lpi_1_dfm_mx0
      = MUX1HOT_s_1_7_2((nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_15_nl),
      Arbiter_8U_Roundrobin_pick_priority_9_sva_1, Arbiter_8U_Roundrobin_pick_priority_11_sva_1,
      (mem_inst_request_xbar_xbar_for_7_lshift_tmp[7]), (mem_inst_request_xbar_xbar_for_1_lshift_tmp[7]),
      (mem_inst_request_xbar_xbar_for_3_lshift_tmp[7]), (mem_inst_request_xbar_xbar_for_5_lshift_tmp[7]),
      {or_dcpl_126 , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_1_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_2_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_3_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_4_nl)
      , (nvhls_leading_ones_3U_nvhls_nvhls_t_3U_nvuint_t_nvhls_nvhls_t_2U_nvuint_t_and_5_nl)});
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_lpi_1_dfm_mx0
      = MUX1HOT_s_1_4_2(Arbiter_8U_Roundrobin_pick_priority_14_sva_1, operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1,
      operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1, operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1,
      {or_dcpl_126 , and_dcpl_339 , and_dcpl_343 , and_dcpl_344});
  assign mem_inst_request_xbar_xbar_for_3_8_operator_3_false_operator_3_false_operator_3_false_or_nl
      = Arbiter_8U_Roundrobin_pick_priority_14_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_12_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_8_operator_4_false_operator_4_false_operator_4_false_or_nl
      = (mem_inst_request_xbar_xbar_for_1_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[7])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[7]);
  assign and_494_nl = or_dcpl_136 & or_dcpl_135 & or_dcpl_134 & or_dcpl_133 & or_dcpl_129
      & or_dcpl_128 & or_dcpl_127;
  assign nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0
      = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_3_8_operator_3_false_operator_3_false_operator_3_false_or_nl),
      (mem_inst_request_xbar_xbar_for_3_8_operator_4_false_operator_4_false_operator_4_false_or_nl),
      and_494_nl);
  assign Arbiter_8U_Roundrobin_pick_priority_9_sva_1 = mem_inst_request_xbar_arbiters_next_7_2_sva
      & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_priority_11_sva_1 = mem_inst_request_xbar_arbiters_next_7_4_sva
      & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[7]);
  assign operator_2_false_operator_2_false_operator_2_false_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_priority_11_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_sva_1;
  assign Arbiter_8U_Roundrobin_pick_priority_10_sva_1 = mem_inst_request_xbar_arbiters_next_7_3_sva
      & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_priority_13_sva_1 = mem_inst_request_xbar_arbiters_next_7_6_sva
      & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_priority_14_sva_1 = mem_inst_request_xbar_arbiters_next_7_7_sva
      & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[7]);
  assign Arbiter_8U_Roundrobin_pick_priority_12_sva_1 = mem_inst_request_xbar_arbiters_next_7_5_sva
      & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[7]);
  assign operator_2_false_1_operator_2_false_1_operator_2_false_1_or_mdf_sva_1 =
      (mem_inst_request_xbar_xbar_for_1_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[7]);
  assign operator_2_false_2_operator_2_false_2_operator_2_false_2_or_mdf_sva_1 =
      (mem_inst_request_xbar_xbar_for_5_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_4_lshift_tmp[7]);
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      = mem_inst_request_xbar_arbiters_next_7_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[7]);
  assign operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1 = Arbiter_8U_Roundrobin_pick_priority_14_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_13_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_sva_1 | Arbiter_8U_Roundrobin_pick_priority_10_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_sva_1 | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1 = ~(mem_inst_request_xbar_xbar_for_3_if_1_mux_28_tmp
      | (~ mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1));
  assign mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1 = ~(mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp
      | (~ mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1));
  assign mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1 = ~(mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp
      | (~ mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1));
  assign mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1 = ~(mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp
      | (~ mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1));
  assign mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1 = ~(mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp
      | (~ mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1));
  assign mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1 = ~(mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp
      | (~ mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1));
  assign mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1 = ~(mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp
      | (~ mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1));
  assign mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1 = ~(mem_inst_request_xbar_xbar_for_3_if_1_mux_tmp
      | (~ mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1));
  assign while_else_while_else_or_10_nl = (while_req_reg_valids_sva_1[7]) | write_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_req_reg_valids_7_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((while_else_while_else_or_10_nl),
      (while_req_reg_valids_sva_1[7]), while_asn_mdf_sva_1);
  assign while_else_while_else_or_11_nl = (while_req_reg_valids_sva_1[6]) | write_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_req_reg_valids_6_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((while_else_while_else_or_11_nl),
      (while_req_reg_valids_sva_1[6]), while_asn_mdf_sva_1);
  assign while_and_21_cse_1 = write_req_PopNB_mioi_return_rsc_z_mxwt & (~ while_asn_mdf_sva_1);
  assign while_else_while_else_or_12_nl = (while_req_reg_valids_sva_1[5]) | write_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_req_reg_valids_5_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((while_else_while_else_or_12_nl),
      (while_req_reg_valids_sva_1[5]), while_asn_mdf_sva_1);
  assign while_else_while_else_or_13_nl = (while_req_reg_valids_sva_1[4]) | write_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_req_reg_valids_4_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((while_else_while_else_or_13_nl),
      (while_req_reg_valids_sva_1[4]), while_asn_mdf_sva_1);
  assign while_else_while_else_or_14_nl = (while_req_reg_valids_sva_1[3]) | write_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_req_reg_valids_3_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((while_else_while_else_or_14_nl),
      (while_req_reg_valids_sva_1[3]), while_asn_mdf_sva_1);
  assign while_else_while_else_or_15_nl = (while_req_reg_valids_sva_1[2]) | write_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_req_reg_valids_2_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((while_else_while_else_or_15_nl),
      (while_req_reg_valids_sva_1[2]), while_asn_mdf_sva_1);
  assign while_else_while_else_or_16_nl = (while_req_reg_valids_sva_1[1]) | write_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_req_reg_valids_1_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((while_else_while_else_or_16_nl),
      (while_req_reg_valids_sva_1[1]), while_asn_mdf_sva_1);
  assign while_else_while_else_or_17_nl = (while_req_reg_valids_sva_1[0]) | write_req_PopNB_mioi_return_rsc_z_mxwt;
  assign while_req_reg_valids_0_lpi_1_dfm_1_mx0 = MUX_s_1_2_2((while_else_while_else_or_17_nl),
      (while_req_reg_valids_sva_1[0]), while_asn_mdf_sva_1);
  assign while_req_reg_type_val_lpi_1_dfm_2 = while_req_reg_type_val_sva_1 | while_and_21_cse_1;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
      = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
      = mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
      = mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
      = mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
      = mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
      = mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
      = mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4;
  assign Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
      = mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5;
  assign mem_inst_load_store_for_4_if_and_tmp_15_sva_1 = mem_inst_load_store_for_4_if_and_stg_1_0_7_sva_1
      & (~ (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[2]));
  assign mem_inst_load_store_for_4_if_and_tmp_7_sva_2 = mem_inst_load_store_for_4_if_and_stg_1_0_sva_1
      & (~ (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[2]));
  assign mem_inst_load_store_for_4_and_41_cse_1 = mem_inst_load_store_for_4_if_and_stg_1_0_1_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_2_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_8_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_3_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_16_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_4_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_24_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_5_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_32_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_6_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_16_m1c_1 = ~(mem_inst_load_store_for_4_and_16_tmp_1
      | mem_inst_load_store_for_4_and_24_tmp_1 | mem_inst_load_store_for_4_and_32_tmp_1);
  assign mem_inst_load_store_for_4_if_and_tmp_14_sva_1 = mem_inst_load_store_for_4_if_and_stg_1_1_7_sva_1
      & (~ (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[2]));
  assign mem_inst_load_store_for_4_if_and_tmp_6_sva_2 = mem_inst_load_store_for_4_if_and_stg_1_1_sva_1
      & (~ (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[2]));
  assign mem_inst_load_store_for_4_and_43_cse_1 = mem_inst_load_store_for_4_if_and_stg_1_1_1_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_1_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_2_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_9_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_3_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_17_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_4_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_25_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_5_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_33_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_6_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_17_m1c_1 = ~(mem_inst_load_store_for_4_and_17_tmp_1
      | mem_inst_load_store_for_4_and_25_tmp_1 | mem_inst_load_store_for_4_and_33_tmp_1);
  assign mem_inst_load_store_for_4_if_and_tmp_13_sva_1 = mem_inst_load_store_for_4_if_and_stg_1_2_7_sva_1
      & (~ (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[2]));
  assign mem_inst_load_store_for_4_if_and_tmp_5_sva_2 = mem_inst_load_store_for_4_if_and_stg_1_2_sva_1
      & (~ (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[2]));
  assign mem_inst_load_store_for_4_and_45_cse_1 = mem_inst_load_store_for_4_if_and_stg_1_2_1_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_2_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_2_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_10_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_3_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_18_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_4_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_26_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_5_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_34_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_6_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_18_m1c_1 = ~(mem_inst_load_store_for_4_and_18_tmp_1
      | mem_inst_load_store_for_4_and_26_tmp_1 | mem_inst_load_store_for_4_and_34_tmp_1);
  assign mem_inst_load_store_for_4_if_and_tmp_12_sva_1 = mem_inst_load_store_for_4_if_and_stg_1_3_7_sva_1
      & (~ (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[2]));
  assign mem_inst_load_store_for_4_if_and_tmp_4_sva_2 = mem_inst_load_store_for_4_if_and_stg_1_3_sva_1
      & (~ (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[2]));
  assign mem_inst_load_store_for_4_and_47_cse_1 = mem_inst_load_store_for_4_if_and_stg_1_3_1_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_3_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_2_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_11_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_3_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_19_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_4_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_27_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_5_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_35_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_6_sva_mx1
      & (~ mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2)
      & mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_19_m1c_1 = ~(mem_inst_load_store_for_4_and_19_tmp_1
      | mem_inst_load_store_for_4_and_27_tmp_1 | mem_inst_load_store_for_4_and_35_tmp_1);
  assign mem_inst_load_store_for_4_if_and_tmp_11_sva_1 = mem_inst_load_store_for_4_if_and_stg_1_0_7_sva_1
      & (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[2]);
  assign mem_inst_load_store_for_4_if_and_tmp_3_sva_2 = mem_inst_load_store_for_4_if_and_stg_1_0_sva_1
      & (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[2]);
  assign mem_inst_load_store_for_4_and_49_cse_1 = mem_inst_load_store_for_4_if_and_stg_1_0_1_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_4_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_2_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_12_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_3_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_20_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_4_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_28_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_5_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_36_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_0_6_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_20_m1c_1 = ~(mem_inst_load_store_for_4_and_20_tmp_1
      | mem_inst_load_store_for_4_and_28_tmp_1 | mem_inst_load_store_for_4_and_36_tmp_1);
  assign mem_inst_load_store_for_4_if_and_tmp_10_sva_1 = mem_inst_load_store_for_4_if_and_stg_1_1_7_sva_1
      & (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[2]);
  assign mem_inst_load_store_for_4_if_and_tmp_2_sva_2 = mem_inst_load_store_for_4_if_and_stg_1_1_sva_1
      & (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[2]);
  assign mem_inst_load_store_for_4_and_51_cse_1 = mem_inst_load_store_for_4_if_and_stg_1_1_1_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_5_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_2_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_13_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_3_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_21_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_4_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_29_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_5_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_37_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_1_6_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_21_m1c_1 = ~(mem_inst_load_store_for_4_and_21_tmp_1
      | mem_inst_load_store_for_4_and_29_tmp_1 | mem_inst_load_store_for_4_and_37_tmp_1);
  assign mem_inst_load_store_for_4_if_and_tmp_9_sva_1 = mem_inst_load_store_for_4_if_and_stg_1_2_7_sva_1
      & (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[2]);
  assign mem_inst_load_store_for_4_if_and_tmp_1_sva_2 = mem_inst_load_store_for_4_if_and_stg_1_2_sva_1
      & (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[2]);
  assign mem_inst_load_store_for_4_and_53_cse_1 = mem_inst_load_store_for_4_if_and_stg_1_2_1_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_6_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_2_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_14_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_3_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_22_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_4_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_30_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_5_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_38_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_2_6_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_22_m1c_1 = ~(mem_inst_load_store_for_4_and_22_tmp_1
      | mem_inst_load_store_for_4_and_30_tmp_1 | mem_inst_load_store_for_4_and_38_tmp_1);
  assign mem_inst_load_store_for_4_if_and_tmp_8_sva_1 = mem_inst_load_store_for_4_if_and_stg_1_3_7_sva_1
      & (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[2]);
  assign mem_inst_load_store_for_4_if_and_tmp_sva_2 = mem_inst_load_store_for_4_if_and_stg_1_3_sva_1
      & (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[2]);
  assign mem_inst_load_store_for_4_and_55_cse_1 = mem_inst_load_store_for_4_if_and_stg_1_3_1_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_7_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_2_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_15_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_3_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_23_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_4_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_31_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_5_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_and_39_tmp_1 = mem_inst_load_store_for_4_if_and_stg_1_3_6_sva_mx1
      & mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx1_2 &
      mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1;
  assign mem_inst_load_store_for_4_mem_inst_load_store_for_4_nor_23_m1c_1 = ~(mem_inst_load_store_for_4_and_23_tmp_1
      | mem_inst_load_store_for_4_and_31_tmp_1 | mem_inst_load_store_for_4_and_39_tmp_1);
  assign mem_inst_load_store_for_4_if_and_stg_1_0_sva_1 = ~((mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[1:0]!=2'b00));
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_3_nl = MUX_v_3_8_2(3'b000, 3'b001,
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_1_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_1_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_1_sva_1});
  assign mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1 = MUX_v_3_2_2(3'b000,
      (mem_inst_request_xbar_xbar_for_3_if_1_mux_3_nl), mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_sva_1 = (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[1:0]==2'b01);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_sva_1 = (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[1:0]==2'b10);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_sva_1 = (mem_inst_request_xbar_run_1_output_data_input_chan_0_lpi_1_dfm_1[1:0]==2'b11);
  assign mem_inst_load_store_for_4_if_or_71_nl = mem_inst_load_store_valid_src_7_lpi_1_dfm_8
      | mem_inst_load_store_for_4_if_and_tmp_8_sva_1;
  assign mem_inst_load_store_valid_src_7_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((mem_inst_load_store_for_4_if_or_71_nl),
      mem_inst_load_store_valid_src_7_lpi_1_dfm_8, or_dcpl_137);
  assign mem_inst_load_store_for_4_if_or_69_nl = mem_inst_load_store_valid_src_6_lpi_1_dfm_8
      | mem_inst_load_store_for_4_if_and_tmp_9_sva_1;
  assign mem_inst_load_store_valid_src_6_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((mem_inst_load_store_for_4_if_or_69_nl),
      mem_inst_load_store_valid_src_6_lpi_1_dfm_8, or_dcpl_137);
  assign mem_inst_load_store_for_4_if_or_67_nl = mem_inst_load_store_valid_src_5_lpi_1_dfm_8
      | mem_inst_load_store_for_4_if_and_tmp_10_sva_1;
  assign mem_inst_load_store_valid_src_5_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((mem_inst_load_store_for_4_if_or_67_nl),
      mem_inst_load_store_valid_src_5_lpi_1_dfm_8, or_dcpl_137);
  assign mem_inst_load_store_for_4_if_or_65_nl = mem_inst_load_store_valid_src_4_lpi_1_dfm_8
      | mem_inst_load_store_for_4_if_and_tmp_11_sva_1;
  assign mem_inst_load_store_valid_src_4_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((mem_inst_load_store_for_4_if_or_65_nl),
      mem_inst_load_store_valid_src_4_lpi_1_dfm_8, or_dcpl_137);
  assign mem_inst_load_store_for_4_if_or_64_nl = mem_inst_load_store_valid_src_3_lpi_1_dfm_8
      | mem_inst_load_store_for_4_if_and_tmp_12_sva_1;
  assign mem_inst_load_store_valid_src_3_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((mem_inst_load_store_for_4_if_or_64_nl),
      mem_inst_load_store_valid_src_3_lpi_1_dfm_8, or_dcpl_137);
  assign mem_inst_load_store_for_4_if_or_66_nl = mem_inst_load_store_valid_src_2_lpi_1_dfm_8
      | mem_inst_load_store_for_4_if_and_tmp_13_sva_1;
  assign mem_inst_load_store_valid_src_2_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((mem_inst_load_store_for_4_if_or_66_nl),
      mem_inst_load_store_valid_src_2_lpi_1_dfm_8, or_dcpl_137);
  assign mem_inst_load_store_for_4_if_or_68_nl = mem_inst_load_store_valid_src_1_lpi_1_dfm_8
      | mem_inst_load_store_for_4_if_and_tmp_14_sva_1;
  assign mem_inst_load_store_valid_src_1_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((mem_inst_load_store_for_4_if_or_68_nl),
      mem_inst_load_store_valid_src_1_lpi_1_dfm_8, or_dcpl_137);
  assign mem_inst_load_store_for_4_if_or_70_nl = mem_inst_load_store_valid_src_0_lpi_1_dfm_8
      | mem_inst_load_store_for_4_if_and_tmp_15_sva_1;
  assign mem_inst_load_store_valid_src_0_lpi_1_dfm_7_mx0 = MUX_s_1_2_2((mem_inst_load_store_for_4_if_or_70_nl),
      mem_inst_load_store_valid_src_0_lpi_1_dfm_8, or_dcpl_137);
  assign mem_inst_load_store_valid_src_7_lpi_1_dfm_8 = (mem_inst_load_store_for_4_if_and_tmp_sva_2
      & mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1) | mem_inst_load_store_for_4_and_55_cse_1
      | mem_inst_load_store_for_4_and_7_tmp_1 | mem_inst_load_store_for_4_and_15_tmp_1
      | mem_inst_load_store_for_4_and_23_tmp_1 | mem_inst_load_store_for_4_and_31_tmp_1
      | mem_inst_load_store_for_4_and_39_tmp_1;
  assign mem_inst_load_store_valid_src_6_lpi_1_dfm_8 = (mem_inst_load_store_for_4_if_and_tmp_1_sva_2
      & mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1) | mem_inst_load_store_for_4_and_53_cse_1
      | mem_inst_load_store_for_4_and_6_tmp_1 | mem_inst_load_store_for_4_and_14_tmp_1
      | mem_inst_load_store_for_4_and_22_tmp_1 | mem_inst_load_store_for_4_and_30_tmp_1
      | mem_inst_load_store_for_4_and_38_tmp_1;
  assign mem_inst_load_store_valid_src_5_lpi_1_dfm_8 = (mem_inst_load_store_for_4_if_and_tmp_2_sva_2
      & mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1) | mem_inst_load_store_for_4_and_51_cse_1
      | mem_inst_load_store_for_4_and_5_tmp_1 | mem_inst_load_store_for_4_and_13_tmp_1
      | mem_inst_load_store_for_4_and_21_tmp_1 | mem_inst_load_store_for_4_and_29_tmp_1
      | mem_inst_load_store_for_4_and_37_tmp_1;
  assign mem_inst_load_store_valid_src_4_lpi_1_dfm_8 = (mem_inst_load_store_for_4_if_and_tmp_3_sva_2
      & mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1) | mem_inst_load_store_for_4_and_49_cse_1
      | mem_inst_load_store_for_4_and_4_tmp_1 | mem_inst_load_store_for_4_and_12_tmp_1
      | mem_inst_load_store_for_4_and_20_tmp_1 | mem_inst_load_store_for_4_and_28_tmp_1
      | mem_inst_load_store_for_4_and_36_tmp_1;
  assign mem_inst_load_store_valid_src_3_lpi_1_dfm_8 = (mem_inst_load_store_for_4_if_and_tmp_4_sva_2
      & mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1) | mem_inst_load_store_for_4_and_47_cse_1
      | mem_inst_load_store_for_4_and_3_tmp_1 | mem_inst_load_store_for_4_and_11_tmp_1
      | mem_inst_load_store_for_4_and_19_tmp_1 | mem_inst_load_store_for_4_and_27_tmp_1
      | mem_inst_load_store_for_4_and_35_tmp_1;
  assign mem_inst_load_store_valid_src_2_lpi_1_dfm_8 = (mem_inst_load_store_for_4_if_and_tmp_5_sva_2
      & mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1) | mem_inst_load_store_for_4_and_45_cse_1
      | mem_inst_load_store_for_4_and_2_tmp_1 | mem_inst_load_store_for_4_and_10_tmp_1
      | mem_inst_load_store_for_4_and_18_tmp_1 | mem_inst_load_store_for_4_and_26_tmp_1
      | mem_inst_load_store_for_4_and_34_tmp_1;
  assign mem_inst_load_store_valid_src_1_lpi_1_dfm_8 = (mem_inst_load_store_for_4_if_and_tmp_6_sva_2
      & mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1) | mem_inst_load_store_for_4_and_43_cse_1
      | mem_inst_load_store_for_4_and_1_tmp_1 | mem_inst_load_store_for_4_and_9_tmp_1
      | mem_inst_load_store_for_4_and_17_tmp_1 | mem_inst_load_store_for_4_and_25_tmp_1
      | mem_inst_load_store_for_4_and_33_tmp_1;
  assign mem_inst_load_store_valid_src_0_lpi_1_dfm_8 = (mem_inst_load_store_for_4_if_and_tmp_7_sva_2
      & mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1) | mem_inst_load_store_for_4_and_41_cse_1
      | mem_inst_load_store_for_4_and_tmp_1 | mem_inst_load_store_for_4_and_8_tmp_1
      | mem_inst_load_store_for_4_and_16_tmp_1 | mem_inst_load_store_for_4_and_24_tmp_1
      | mem_inst_load_store_for_4_and_32_tmp_1;
  assign mem_inst_load_store_for_4_if_and_stg_1_0_7_sva_1 = ~((mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[1:0]!=2'b00));
  assign mem_inst_request_xbar_xbar_for_3_if_1_mux_31_nl = MUX_v_3_8_2(3'b000, 3'b001,
      3'b010, 3'b011, 3'b100, 3'b101, 3'b110, 3'b111, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_sva_1});
  assign mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2 = MUX_v_3_2_2(3'b000,
      (mem_inst_request_xbar_xbar_for_3_if_1_mux_31_nl), mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1);
  assign mem_inst_load_store_for_4_if_and_stg_1_1_7_sva_1 = (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[1:0]==2'b01);
  assign mem_inst_load_store_for_4_if_and_stg_1_2_7_sva_1 = (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[1:0]==2'b10);
  assign mem_inst_load_store_for_4_if_and_stg_1_3_7_sva_1 = (mem_inst_request_xbar_run_1_output_data_input_chan_7_lpi_1_dfm_2[1:0]==2'b11);
  assign Arbiter_8U_Roundrobin_pick_if_1_not_64 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1);
  assign and_dcpl = while_stage_0_5 & while_asn_mdf_sva_st_1_3;
  assign and_dcpl_1 = while_stage_0_4 & while_lor_lpi_1_dfm_st_1;
  assign or_dcpl_1 = while_asn_mdf_sva_st_1_2 | (~ while_stage_0_3) | (~ while_if_1_while_if_1_or_tmp);
  assign nor_tmp_1 = while_asn_mdf_sva_st_1_2 & while_stage_0_4;
  assign and_685_cse = while_if_1_while_if_1_or_tmp & while_stage_0_3;
  assign and_tmp = Arbiter_8U_Roundrobin_pick_unequal_tmp_8 & (mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2
      | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1);
  assign and_tmp_1 = Arbiter_8U_Roundrobin_pick_unequal_tmp_9 & (mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0);
  assign and_tmp_2 = Arbiter_8U_Roundrobin_pick_unequal_tmp_10 & (mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2
      | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1);
  assign and_tmp_3 = (mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7)
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_11;
  assign and_tmp_4 = (mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4)
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_12;
  assign and_tmp_5 = (mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7)
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_13;
  assign and_tmp_6 = (mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7)
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_14;
  assign and_tmp_7 = (mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_5
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_4
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_2
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_0
      | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_3)
      & Arbiter_8U_Roundrobin_pick_unequal_tmp_15;
  assign or_dcpl_11 = ~(while_lor_lpi_1_dfm_2 & while_stage_0_5);
  assign or_dcpl_12 = ~(while_stage_0_3 & while_if_1_while_if_1_or_tmp);
  assign and_dcpl_122 = ~((mem_inst_request_xbar_xbar_for_1_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[0])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[0]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[0]));
  assign and_dcpl_131 = ~((mem_inst_request_xbar_xbar_for_7_lshift_tmp[1]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[1]));
  assign and_dcpl_134 = ~((mem_inst_request_xbar_xbar_for_1_lshift_tmp[2]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[2]));
  assign and_dcpl_144 = ~((mem_inst_request_xbar_xbar_for_7_lshift_tmp[3]) | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[3]));
  assign and_dcpl_148 = ~((mem_inst_request_xbar_xbar_for_1_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[4]));
  assign and_dcpl_151 = ~((mem_inst_request_xbar_xbar_for_6_lshift_tmp[4]) | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[4]));
  assign and_dcpl_157 = ~((mem_inst_request_xbar_xbar_for_8_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[5])
      | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[5]) | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[5]));
  assign and_dcpl_167 = ~((mem_inst_request_xbar_xbar_for_1_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[6])
      | (mem_inst_request_xbar_xbar_for_6_lshift_tmp[6]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[6]));
  assign and_dcpl_171 = ~((mem_inst_request_xbar_xbar_for_6_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_1_lshift_tmp[7])
      | (mem_inst_request_xbar_xbar_for_7_lshift_tmp[7]) | (mem_inst_request_xbar_xbar_for_8_lshift_tmp[7]));
  assign or_dcpl_24 = (~ and_tmp_1) | mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp;
  assign or_dcpl_27 = (~ and_tmp_2) | mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp;
  assign or_dcpl_30 = (~ and_tmp_3) | mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp;
  assign or_dcpl_33 = (~ and_tmp_4) | mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp;
  assign or_dcpl_36 = (~ and_tmp_5) | mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp;
  assign or_dcpl_39 = (~ and_tmp_6) | mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp;
  assign or_dcpl_40 = while_asn_mdf_sva_1 | (~ write_req_PopNB_mioi_return_rsc_z_mxwt);
  assign or_dcpl_41 = Arbiter_8U_Roundrobin_pick_priority_12_1_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_1_sva_1;
  assign or_dcpl_42 = or_dcpl_41 | Arbiter_8U_Roundrobin_pick_priority_14_1_sva_1;
  assign or_dcpl_43 = ~(mem_inst_request_xbar_arbiters_next_0_7_sva & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[0]));
  assign or_dcpl_44 = ~(mem_inst_request_xbar_arbiters_next_0_6_sva & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[0]));
  assign or_dcpl_45 = ~(mem_inst_request_xbar_arbiters_next_0_5_sva & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[0]));
  assign or_dcpl_47 = mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | Arbiter_8U_Roundrobin_pick_priority_9_1_sva_1;
  assign and_dcpl_185 = (or_dcpl_47 | Arbiter_8U_Roundrobin_pick_priority_10_1_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_1_sva_1) & or_dcpl_45 & or_dcpl_44
      & or_dcpl_43;
  assign or_dcpl_49 = ~(mem_inst_request_xbar_arbiters_next_0_4_sva & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[0]));
  assign or_dcpl_50 = ~(mem_inst_request_xbar_arbiters_next_0_3_sva & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[0]));
  assign or_dcpl_51 = ~(mem_inst_request_xbar_arbiters_next_0_2_sva & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[0]));
  assign or_dcpl_52 = ~((mem_inst_request_xbar_xbar_for_2_lshift_tmp[0]) & mem_inst_request_xbar_arbiters_next_0_1_sva);
  assign mux_1_nl = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_1_lshift_tmp[0]),
      (~ mem_inst_request_xbar_arbiters_next_0_5_sva), mem_inst_request_xbar_xbar_for_6_lshift_tmp[0]);
  assign nor_45_nl = ~(mem_inst_request_xbar_arbiters_next_0_6_sva | Arbiter_8U_Roundrobin_pick_priority_12_1_sva_1);
  assign mux_2_nl = MUX_s_1_2_2((mux_1_nl), (nor_45_nl), mem_inst_request_xbar_xbar_for_7_lshift_tmp[0]);
  assign nor_46_nl = ~(mem_inst_request_xbar_arbiters_next_0_7_sva | or_dcpl_41);
  assign mux_3_nl = MUX_s_1_2_2((mux_2_nl), (nor_46_nl), mem_inst_request_xbar_xbar_for_8_lshift_tmp[0]);
  assign and_dcpl_189 = (mux_3_nl) & or_dcpl_52 & or_dcpl_51 & or_dcpl_50 & or_dcpl_49;
  assign nor_38_nl = ~(mem_inst_request_xbar_arbiters_next_0_1_sva | (~ (mem_inst_request_xbar_xbar_for_2_lshift_tmp[0])));
  assign nor_39_nl = ~(mem_inst_request_xbar_arbiters_next_0_2_sva | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_priority_and_5_cse);
  assign mux_4_nl = MUX_s_1_2_2((nor_38_nl), (nor_39_nl), mem_inst_request_xbar_xbar_for_3_lshift_tmp[0]);
  assign nor_40_nl = ~(mem_inst_request_xbar_arbiters_next_0_3_sva | or_dcpl_47);
  assign mux_5_nl = MUX_s_1_2_2((mux_4_nl), (nor_40_nl), mem_inst_request_xbar_xbar_for_4_lshift_tmp[0]);
  assign nor_41_nl = ~(mem_inst_request_xbar_arbiters_next_0_4_sva | Arbiter_8U_Roundrobin_pick_priority_10_1_sva_1
      | or_dcpl_47);
  assign mux_6_nl = MUX_s_1_2_2((mux_5_nl), (nor_41_nl), mem_inst_request_xbar_xbar_for_5_lshift_tmp[0]);
  assign and_dcpl_190 = (mux_6_nl) & and_dcpl_122;
  assign or_dcpl_53 = Arbiter_8U_Roundrobin_pick_priority_13_2_sva_1 | Arbiter_8U_Roundrobin_pick_priority_14_2_sva_1;
  assign or_dcpl_54 = or_dcpl_53 | Arbiter_8U_Roundrobin_pick_priority_12_2_sva_1;
  assign or_dcpl_55 = ~(mem_inst_request_xbar_arbiters_next_1_5_sva & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[1]));
  assign or_dcpl_56 = ~(mem_inst_request_xbar_arbiters_next_1_7_sva & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[1]));
  assign or_dcpl_57 = ~((mem_inst_request_xbar_xbar_for_7_lshift_tmp[1]) & mem_inst_request_xbar_arbiters_next_1_6_sva);
  assign and_dcpl_206 = (operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1
      | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | Arbiter_8U_Roundrobin_pick_priority_9_2_sva_1) & or_dcpl_57 & or_dcpl_56
      & or_dcpl_55;
  assign or_dcpl_61 = ~(mem_inst_request_xbar_arbiters_next_1_2_sva & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[1]));
  assign or_dcpl_62 = ~(mem_inst_request_xbar_arbiters_next_1_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[1]));
  assign or_dcpl_63 = ~(mem_inst_request_xbar_arbiters_next_1_3_sva & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[1]));
  assign or_dcpl_64 = ~((mem_inst_request_xbar_xbar_for_5_lshift_tmp[1]) & mem_inst_request_xbar_arbiters_next_1_4_sva);
  assign or_171_nl = mem_inst_request_xbar_arbiters_next_1_6_sva | (~ (mem_inst_request_xbar_xbar_for_7_lshift_tmp[1]));
  assign or_170_nl = mem_inst_request_xbar_arbiters_next_1_7_sva | Arbiter_8U_Roundrobin_pick_priority_13_2_sva_1;
  assign mux_7_nl = MUX_s_1_2_2((or_171_nl), (or_170_nl), mem_inst_request_xbar_xbar_for_8_lshift_tmp[1]);
  assign mux_8_nl = MUX_s_1_2_2((mux_7_nl), or_dcpl_53, mem_inst_request_xbar_xbar_for_1_lshift_tmp[1]);
  assign or_169_nl = mem_inst_request_xbar_arbiters_next_1_5_sva | or_dcpl_53;
  assign mux_9_nl = MUX_s_1_2_2((mux_8_nl), (or_169_nl), mem_inst_request_xbar_xbar_for_6_lshift_tmp[1]);
  assign and_dcpl_210 = (~ (mux_9_nl)) & or_dcpl_64 & or_dcpl_63 & or_dcpl_62 & or_dcpl_61;
  assign nor_34_nl = ~(mem_inst_request_xbar_arbiters_next_1_4_sva | (~ (mem_inst_request_xbar_xbar_for_5_lshift_tmp[1])));
  assign nor_35_nl = ~(mem_inst_request_xbar_arbiters_next_1_3_sva | Arbiter_8U_Roundrobin_pick_priority_11_2_sva_1);
  assign mux_10_nl = MUX_s_1_2_2((nor_34_nl), (nor_35_nl), mem_inst_request_xbar_xbar_for_4_lshift_tmp[1]);
  assign nor_36_nl = ~(mem_inst_request_xbar_arbiters_next_1_1_sva | operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1);
  assign mux_11_nl = MUX_s_1_2_2((mux_10_nl), (nor_36_nl), mem_inst_request_xbar_xbar_for_2_lshift_tmp[1]);
  assign nor_37_nl = ~(mem_inst_request_xbar_arbiters_next_1_2_sva | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | operator_2_false_operator_2_false_operator_2_false_or_mdf_2_sva_1);
  assign mux_12_nl = MUX_s_1_2_2((mux_11_nl), (nor_37_nl), mem_inst_request_xbar_xbar_for_3_lshift_tmp[1]);
  assign and_dcpl_213 = (mux_12_nl) & and_dcpl_131 & (~ (mem_inst_request_xbar_xbar_for_1_lshift_tmp[1]))
      & (~ (mem_inst_request_xbar_xbar_for_6_lshift_tmp[1]));
  assign or_dcpl_65 = Arbiter_8U_Roundrobin_pick_priority_12_3_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_3_sva_1;
  assign or_dcpl_66 = or_dcpl_65 | Arbiter_8U_Roundrobin_pick_priority_14_3_sva_1;
  assign or_dcpl_67 = ~(mem_inst_request_xbar_arbiters_next_2_7_sva & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[2]));
  assign or_dcpl_68 = ~(mem_inst_request_xbar_arbiters_next_2_6_sva & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[2]));
  assign or_dcpl_69 = ~((mem_inst_request_xbar_xbar_for_6_lshift_tmp[2]) & mem_inst_request_xbar_arbiters_next_2_5_sva);
  assign and_dcpl_229 = (operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_9_3_sva_1 | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_priority_and_5_cse)
      & or_dcpl_69 & or_dcpl_68 & or_dcpl_67;
  assign or_dcpl_73 = ~(mem_inst_request_xbar_arbiters_next_2_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[2]));
  assign or_dcpl_74 = ~(mem_inst_request_xbar_arbiters_next_2_2_sva & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[2]));
  assign or_dcpl_75 = ~(mem_inst_request_xbar_arbiters_next_2_3_sva & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[2]));
  assign or_dcpl_76 = ~((mem_inst_request_xbar_xbar_for_5_lshift_tmp[2]) & mem_inst_request_xbar_arbiters_next_2_4_sva);
  assign or_191_nl = mem_inst_request_xbar_arbiters_next_2_5_sva | (~ (mem_inst_request_xbar_xbar_for_6_lshift_tmp[2]));
  assign or_190_nl = mem_inst_request_xbar_arbiters_next_2_6_sva | Arbiter_8U_Roundrobin_pick_priority_12_3_sva_1;
  assign mux_13_nl = MUX_s_1_2_2((or_191_nl), (or_190_nl), mem_inst_request_xbar_xbar_for_7_lshift_tmp[2]);
  assign mux_14_nl = MUX_s_1_2_2((mux_13_nl), or_dcpl_65, mem_inst_request_xbar_xbar_for_1_lshift_tmp[2]);
  assign or_189_nl = mem_inst_request_xbar_arbiters_next_2_7_sva | or_dcpl_65;
  assign mux_15_nl = MUX_s_1_2_2((mux_14_nl), (or_189_nl), mem_inst_request_xbar_xbar_for_8_lshift_tmp[2]);
  assign and_dcpl_233 = (~ (mux_15_nl)) & or_dcpl_76 & or_dcpl_75 & or_dcpl_74 &
      or_dcpl_73;
  assign nor_30_nl = ~(mem_inst_request_xbar_arbiters_next_2_4_sva | (~ (mem_inst_request_xbar_xbar_for_5_lshift_tmp[2])));
  assign nor_31_nl = ~(mem_inst_request_xbar_arbiters_next_2_3_sva | Arbiter_8U_Roundrobin_pick_priority_11_3_sva_1);
  assign mux_16_nl = MUX_s_1_2_2((nor_30_nl), (nor_31_nl), mem_inst_request_xbar_xbar_for_4_lshift_tmp[2]);
  assign nor_32_nl = ~(mem_inst_request_xbar_arbiters_next_2_2_sva | operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1);
  assign mux_17_nl = MUX_s_1_2_2((mux_16_nl), (nor_32_nl), mem_inst_request_xbar_xbar_for_3_lshift_tmp[2]);
  assign nor_33_nl = ~(mem_inst_request_xbar_arbiters_next_2_1_sva | Arbiter_8U_Roundrobin_pick_priority_9_3_sva_1
      | operator_2_false_operator_2_false_operator_2_false_or_mdf_3_sva_1);
  assign mux_18_nl = MUX_s_1_2_2((mux_17_nl), (nor_33_nl), mem_inst_request_xbar_xbar_for_2_lshift_tmp[2]);
  assign and_dcpl_236 = (mux_18_nl) & (~ (mem_inst_request_xbar_xbar_for_6_lshift_tmp[2]))
      & (~ (mem_inst_request_xbar_xbar_for_7_lshift_tmp[2])) & and_dcpl_134;
  assign or_dcpl_77 = Arbiter_8U_Roundrobin_pick_priority_13_4_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_4_sva_1;
  assign or_dcpl_78 = or_dcpl_77 | Arbiter_8U_Roundrobin_pick_priority_14_4_sva_1;
  assign or_dcpl_79 = ~(mem_inst_request_xbar_arbiters_next_3_7_sva & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[3]));
  assign or_dcpl_80 = ~(mem_inst_request_xbar_arbiters_next_3_5_sva & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[3]));
  assign or_dcpl_81 = ~((mem_inst_request_xbar_xbar_for_7_lshift_tmp[3]) & mem_inst_request_xbar_arbiters_next_3_6_sva);
  assign and_dcpl_252 = (operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1
      | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | Arbiter_8U_Roundrobin_pick_priority_9_4_sva_1) & or_dcpl_81 & or_dcpl_80
      & or_dcpl_79;
  assign or_dcpl_85 = ~(mem_inst_request_xbar_arbiters_next_3_2_sva & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[3]));
  assign or_dcpl_86 = ~(mem_inst_request_xbar_arbiters_next_3_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[3]));
  assign or_dcpl_87 = ~(mem_inst_request_xbar_arbiters_next_3_3_sva & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[3]));
  assign or_dcpl_88 = ~((mem_inst_request_xbar_xbar_for_5_lshift_tmp[3]) & mem_inst_request_xbar_arbiters_next_3_4_sva);
  assign or_211_nl = mem_inst_request_xbar_arbiters_next_3_6_sva | (~ (mem_inst_request_xbar_xbar_for_7_lshift_tmp[3]));
  assign or_210_nl = mem_inst_request_xbar_arbiters_next_3_5_sva | Arbiter_8U_Roundrobin_pick_priority_13_4_sva_1;
  assign mux_19_nl = MUX_s_1_2_2((or_211_nl), (or_210_nl), mem_inst_request_xbar_xbar_for_6_lshift_tmp[3]);
  assign or_209_nl = mem_inst_request_xbar_arbiters_next_3_7_sva | or_dcpl_77;
  assign mux_20_nl = MUX_s_1_2_2((mux_19_nl), (or_209_nl), mem_inst_request_xbar_xbar_for_8_lshift_tmp[3]);
  assign mux_21_nl = MUX_s_1_2_2((mux_20_nl), or_dcpl_78, mem_inst_request_xbar_xbar_for_1_lshift_tmp[3]);
  assign and_dcpl_256 = (~ (mux_21_nl)) & or_dcpl_88 & or_dcpl_87 & or_dcpl_86 &
      or_dcpl_85;
  assign nor_26_nl = ~(mem_inst_request_xbar_arbiters_next_3_4_sva | (~ (mem_inst_request_xbar_xbar_for_5_lshift_tmp[3])));
  assign nor_27_nl = ~(mem_inst_request_xbar_arbiters_next_3_3_sva | Arbiter_8U_Roundrobin_pick_priority_11_4_sva_1);
  assign mux_22_nl = MUX_s_1_2_2((nor_26_nl), (nor_27_nl), mem_inst_request_xbar_xbar_for_4_lshift_tmp[3]);
  assign nor_28_nl = ~(mem_inst_request_xbar_arbiters_next_3_1_sva | operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1);
  assign mux_23_nl = MUX_s_1_2_2((mux_22_nl), (nor_28_nl), mem_inst_request_xbar_xbar_for_2_lshift_tmp[3]);
  assign nor_29_nl = ~(mem_inst_request_xbar_arbiters_next_3_2_sva | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | operator_2_false_operator_2_false_operator_2_false_or_mdf_4_sva_1);
  assign mux_24_nl = MUX_s_1_2_2((mux_23_nl), (nor_29_nl), mem_inst_request_xbar_xbar_for_3_lshift_tmp[3]);
  assign and_dcpl_259 = (mux_24_nl) & and_dcpl_144 & (~ (mem_inst_request_xbar_xbar_for_8_lshift_tmp[3]))
      & (~ (mem_inst_request_xbar_xbar_for_1_lshift_tmp[3]));
  assign or_dcpl_89 = Arbiter_8U_Roundrobin_pick_priority_12_5_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_5_sva_1;
  assign or_dcpl_90 = or_dcpl_89 | Arbiter_8U_Roundrobin_pick_priority_14_5_sva_1;
  assign or_dcpl_91 = ~(mem_inst_request_xbar_arbiters_next_4_7_sva & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[4]));
  assign or_dcpl_92 = ~(mem_inst_request_xbar_arbiters_next_4_6_sva & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[4]));
  assign or_dcpl_93 = ~((mem_inst_request_xbar_xbar_for_6_lshift_tmp[4]) & mem_inst_request_xbar_arbiters_next_4_5_sva);
  assign and_dcpl_275 = (operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1
      | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | Arbiter_8U_Roundrobin_pick_priority_9_5_sva_1) & or_dcpl_93 & or_dcpl_92
      & or_dcpl_91;
  assign or_dcpl_97 = ~(mem_inst_request_xbar_arbiters_next_4_2_sva & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[4]));
  assign or_dcpl_98 = ~(mem_inst_request_xbar_arbiters_next_4_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[4]));
  assign or_dcpl_99 = ~(mem_inst_request_xbar_arbiters_next_4_4_sva & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[4]));
  assign or_dcpl_100 = ~((mem_inst_request_xbar_xbar_for_4_lshift_tmp[4]) & mem_inst_request_xbar_arbiters_next_4_3_sva);
  assign or_231_nl = mem_inst_request_xbar_arbiters_next_4_5_sva | (~ (mem_inst_request_xbar_xbar_for_6_lshift_tmp[4]));
  assign or_230_nl = mem_inst_request_xbar_arbiters_next_4_6_sva | Arbiter_8U_Roundrobin_pick_priority_12_5_sva_1;
  assign mux_25_nl = MUX_s_1_2_2((or_231_nl), (or_230_nl), mem_inst_request_xbar_xbar_for_7_lshift_tmp[4]);
  assign mux_26_nl = MUX_s_1_2_2((mux_25_nl), or_dcpl_89, mem_inst_request_xbar_xbar_for_1_lshift_tmp[4]);
  assign or_229_nl = mem_inst_request_xbar_arbiters_next_4_7_sva | or_dcpl_89;
  assign mux_27_nl = MUX_s_1_2_2((mux_26_nl), (or_229_nl), mem_inst_request_xbar_xbar_for_8_lshift_tmp[4]);
  assign and_dcpl_279 = (~ (mux_27_nl)) & or_dcpl_100 & or_dcpl_99 & or_dcpl_98 &
      or_dcpl_97;
  assign nor_22_nl = ~(mem_inst_request_xbar_arbiters_next_4_3_sva | (~ (mem_inst_request_xbar_xbar_for_4_lshift_tmp[4])));
  assign nor_23_nl = ~(mem_inst_request_xbar_arbiters_next_4_4_sva | Arbiter_8U_Roundrobin_pick_priority_10_5_sva_1);
  assign mux_28_nl = MUX_s_1_2_2((nor_22_nl), (nor_23_nl), mem_inst_request_xbar_xbar_for_5_lshift_tmp[4]);
  assign nor_24_nl = ~(mem_inst_request_xbar_arbiters_next_4_1_sva | operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1);
  assign mux_29_nl = MUX_s_1_2_2((mux_28_nl), (nor_24_nl), mem_inst_request_xbar_xbar_for_2_lshift_tmp[4]);
  assign nor_25_nl = ~(mem_inst_request_xbar_arbiters_next_4_2_sva | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | operator_2_false_operator_2_false_operator_2_false_or_mdf_5_sva_1);
  assign mux_30_nl = MUX_s_1_2_2((mux_29_nl), (nor_25_nl), mem_inst_request_xbar_xbar_for_3_lshift_tmp[4]);
  assign and_dcpl_281 = (mux_30_nl) & and_dcpl_151 & and_dcpl_148;
  assign or_dcpl_101 = Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_6_sva_1;
  assign or_dcpl_102 = or_dcpl_101 | Arbiter_8U_Roundrobin_pick_priority_13_6_sva_1;
  assign or_dcpl_103 = ~(mem_inst_request_xbar_arbiters_next_5_6_sva & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[5]));
  assign or_dcpl_104 = ~(mem_inst_request_xbar_arbiters_next_5_5_sva & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[5]));
  assign or_dcpl_105 = ~(mem_inst_request_xbar_arbiters_next_5_7_sva & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[5]));
  assign or_dcpl_107 = mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | Arbiter_8U_Roundrobin_pick_priority_9_6_sva_1;
  assign and_dcpl_297 = (or_dcpl_107 | Arbiter_8U_Roundrobin_pick_priority_10_6_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_11_6_sva_1) & or_dcpl_105 & or_dcpl_104
      & or_dcpl_103;
  assign or_dcpl_109 = ~(mem_inst_request_xbar_arbiters_next_5_4_sva & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[5]));
  assign or_dcpl_110 = ~(mem_inst_request_xbar_arbiters_next_5_3_sva & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[5]));
  assign or_dcpl_111 = ~(mem_inst_request_xbar_arbiters_next_5_2_sva & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[5]));
  assign or_dcpl_112 = ~((mem_inst_request_xbar_xbar_for_2_lshift_tmp[5]) & mem_inst_request_xbar_arbiters_next_5_1_sva);
  assign or_251_nl = (~ (mem_inst_request_xbar_xbar_for_8_lshift_tmp[5])) | mem_inst_request_xbar_arbiters_next_5_7_sva;
  assign mux_31_nl = MUX_s_1_2_2((or_251_nl), Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1,
      mem_inst_request_xbar_xbar_for_1_lshift_tmp[5]);
  assign or_250_nl = mem_inst_request_xbar_arbiters_next_5_5_sva | Arbiter_8U_Roundrobin_pick_priority_14_6_sva_1;
  assign mux_32_nl = MUX_s_1_2_2((mux_31_nl), (or_250_nl), mem_inst_request_xbar_xbar_for_6_lshift_tmp[5]);
  assign or_249_nl = mem_inst_request_xbar_arbiters_next_5_6_sva | or_dcpl_101;
  assign mux_33_nl = MUX_s_1_2_2((mux_32_nl), (or_249_nl), mem_inst_request_xbar_xbar_for_7_lshift_tmp[5]);
  assign and_dcpl_301 = (~ (mux_33_nl)) & or_dcpl_112 & or_dcpl_111 & or_dcpl_110
      & or_dcpl_109;
  assign nor_18_nl = ~(mem_inst_request_xbar_arbiters_next_5_1_sva | (~ (mem_inst_request_xbar_xbar_for_2_lshift_tmp[5])));
  assign nor_19_nl = ~(mem_inst_request_xbar_arbiters_next_5_2_sva | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_priority_and_5_cse);
  assign mux_34_nl = MUX_s_1_2_2((nor_18_nl), (nor_19_nl), mem_inst_request_xbar_xbar_for_3_lshift_tmp[5]);
  assign nor_20_nl = ~(mem_inst_request_xbar_arbiters_next_5_3_sva | or_dcpl_107);
  assign mux_35_nl = MUX_s_1_2_2((mux_34_nl), (nor_20_nl), mem_inst_request_xbar_xbar_for_4_lshift_tmp[5]);
  assign nor_21_nl = ~(mem_inst_request_xbar_arbiters_next_5_4_sva | Arbiter_8U_Roundrobin_pick_priority_10_6_sva_1
      | or_dcpl_107);
  assign mux_36_nl = MUX_s_1_2_2((mux_35_nl), (nor_21_nl), mem_inst_request_xbar_xbar_for_5_lshift_tmp[5]);
  assign and_dcpl_302 = (mux_36_nl) & and_dcpl_157;
  assign or_dcpl_113 = Arbiter_8U_Roundrobin_pick_priority_13_7_sva_1 | Arbiter_8U_Roundrobin_pick_priority_12_7_sva_1;
  assign or_dcpl_114 = or_dcpl_113 | Arbiter_8U_Roundrobin_pick_priority_14_7_sva_1;
  assign or_dcpl_115 = ~(mem_inst_request_xbar_arbiters_next_6_7_sva & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[6]));
  assign or_dcpl_116 = ~(mem_inst_request_xbar_arbiters_next_6_5_sva & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[6]));
  assign or_dcpl_117 = ~(mem_inst_request_xbar_arbiters_next_6_6_sva & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[6]));
  assign and_dcpl_318 = (operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1
      | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | Arbiter_8U_Roundrobin_pick_priority_9_7_sva_1) & or_dcpl_117 & or_dcpl_116
      & or_dcpl_115;
  assign or_dcpl_121 = ~(mem_inst_request_xbar_arbiters_next_6_2_sva & (mem_inst_request_xbar_xbar_for_3_lshift_tmp[6]));
  assign or_dcpl_122 = ~(mem_inst_request_xbar_arbiters_next_6_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[6]));
  assign or_dcpl_123 = ~(mem_inst_request_xbar_arbiters_next_6_4_sva & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[6]));
  assign or_dcpl_124 = ~(mem_inst_request_xbar_arbiters_next_6_3_sva & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[6]));
  assign mux_37_nl = MUX_s_1_2_2((mem_inst_request_xbar_xbar_for_1_lshift_tmp[6]),
      (~ mem_inst_request_xbar_arbiters_next_6_6_sva), mem_inst_request_xbar_xbar_for_7_lshift_tmp[6]);
  assign nor_nl = ~(mem_inst_request_xbar_arbiters_next_6_5_sva | Arbiter_8U_Roundrobin_pick_priority_13_7_sva_1);
  assign mux_38_nl = MUX_s_1_2_2((mux_37_nl), (nor_nl), mem_inst_request_xbar_xbar_for_6_lshift_tmp[6]);
  assign nor_42_nl = ~(mem_inst_request_xbar_arbiters_next_6_7_sva | or_dcpl_113);
  assign mux_39_nl = MUX_s_1_2_2((mux_38_nl), (nor_42_nl), mem_inst_request_xbar_xbar_for_8_lshift_tmp[6]);
  assign and_dcpl_322 = (mux_39_nl) & or_dcpl_124 & or_dcpl_123 & or_dcpl_122 & or_dcpl_121;
  assign nor_14_nl = ~((~ (mem_inst_request_xbar_xbar_for_4_lshift_tmp[6])) | mem_inst_request_xbar_arbiters_next_6_3_sva);
  assign nor_15_nl = ~(mem_inst_request_xbar_arbiters_next_6_4_sva | Arbiter_8U_Roundrobin_pick_priority_10_7_sva_1);
  assign mux_40_nl = MUX_s_1_2_2((nor_14_nl), (nor_15_nl), mem_inst_request_xbar_xbar_for_5_lshift_tmp[6]);
  assign nor_16_nl = ~(mem_inst_request_xbar_arbiters_next_6_1_sva | operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1);
  assign mux_41_nl = MUX_s_1_2_2((mux_40_nl), (nor_16_nl), mem_inst_request_xbar_xbar_for_2_lshift_tmp[6]);
  assign nor_17_nl = ~(mem_inst_request_xbar_arbiters_next_6_2_sva | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_priority_and_5_cse
      | operator_2_false_operator_2_false_operator_2_false_or_mdf_7_sva_1);
  assign mux_42_nl = MUX_s_1_2_2((mux_41_nl), (nor_17_nl), mem_inst_request_xbar_xbar_for_3_lshift_tmp[6]);
  assign and_dcpl_323 = (mux_42_nl) & and_dcpl_167;
  assign or_dcpl_125 = Arbiter_8U_Roundrobin_pick_priority_12_sva_1 | Arbiter_8U_Roundrobin_pick_priority_13_sva_1;
  assign or_dcpl_126 = or_dcpl_125 | Arbiter_8U_Roundrobin_pick_priority_14_sva_1;
  assign or_dcpl_127 = ~(mem_inst_request_xbar_arbiters_next_7_7_sva & (mem_inst_request_xbar_xbar_for_8_lshift_tmp[7]));
  assign or_dcpl_128 = ~(mem_inst_request_xbar_arbiters_next_7_6_sva & (mem_inst_request_xbar_xbar_for_7_lshift_tmp[7]));
  assign or_dcpl_129 = ~(mem_inst_request_xbar_arbiters_next_7_5_sva & (mem_inst_request_xbar_xbar_for_6_lshift_tmp[7]));
  assign or_dcpl_131 = Arbiter_8U_Roundrobin_pick_priority_9_sva_1 | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_priority_and_5_cse;
  assign and_dcpl_339 = (or_dcpl_131 | Arbiter_8U_Roundrobin_pick_priority_11_sva_1
      | Arbiter_8U_Roundrobin_pick_priority_10_sva_1) & or_dcpl_129 & or_dcpl_128
      & or_dcpl_127;
  assign or_dcpl_133 = ~(mem_inst_request_xbar_arbiters_next_7_3_sva & (mem_inst_request_xbar_xbar_for_4_lshift_tmp[7]));
  assign or_dcpl_134 = ~(mem_inst_request_xbar_arbiters_next_7_4_sva & (mem_inst_request_xbar_xbar_for_5_lshift_tmp[7]));
  assign or_dcpl_135 = ~(mem_inst_request_xbar_arbiters_next_7_1_sva & (mem_inst_request_xbar_xbar_for_2_lshift_tmp[7]));
  assign or_dcpl_136 = ~((mem_inst_request_xbar_xbar_for_3_lshift_tmp[7]) & mem_inst_request_xbar_arbiters_next_7_2_sva);
  assign or_290_nl = (~ (mem_inst_request_xbar_xbar_for_6_lshift_tmp[7])) | mem_inst_request_xbar_arbiters_next_7_5_sva;
  assign mux_43_nl = MUX_s_1_2_2((or_290_nl), Arbiter_8U_Roundrobin_pick_priority_12_sva_1,
      mem_inst_request_xbar_xbar_for_1_lshift_tmp[7]);
  assign or_289_nl = mem_inst_request_xbar_arbiters_next_7_6_sva | Arbiter_8U_Roundrobin_pick_priority_12_sva_1;
  assign mux_44_nl = MUX_s_1_2_2((mux_43_nl), (or_289_nl), mem_inst_request_xbar_xbar_for_7_lshift_tmp[7]);
  assign or_288_nl = mem_inst_request_xbar_arbiters_next_7_7_sva | or_dcpl_125;
  assign mux_45_nl = MUX_s_1_2_2((mux_44_nl), (or_288_nl), mem_inst_request_xbar_xbar_for_8_lshift_tmp[7]);
  assign and_dcpl_343 = (~ (mux_45_nl)) & or_dcpl_136 & or_dcpl_135 & or_dcpl_134
      & or_dcpl_133;
  assign nor_10_nl = ~(mem_inst_request_xbar_arbiters_next_7_2_sva | (~ (mem_inst_request_xbar_xbar_for_3_lshift_tmp[7])));
  assign nor_11_nl = ~(mem_inst_request_xbar_arbiters_next_7_1_sva | Arbiter_8U_Roundrobin_pick_priority_9_sva_1);
  assign mux_46_nl = MUX_s_1_2_2((nor_10_nl), (nor_11_nl), mem_inst_request_xbar_xbar_for_2_lshift_tmp[7]);
  assign nor_12_nl = ~(mem_inst_request_xbar_arbiters_next_7_4_sva | or_dcpl_131);
  assign mux_47_nl = MUX_s_1_2_2((mux_46_nl), (nor_12_nl), mem_inst_request_xbar_xbar_for_5_lshift_tmp[7]);
  assign nor_13_nl = ~(mem_inst_request_xbar_arbiters_next_7_3_sva | Arbiter_8U_Roundrobin_pick_priority_11_sva_1
      | or_dcpl_131);
  assign mux_48_nl = MUX_s_1_2_2((mux_47_nl), (nor_13_nl), mem_inst_request_xbar_xbar_for_4_lshift_tmp[7]);
  assign and_dcpl_344 = (mux_48_nl) & and_dcpl_171;
  assign or_dcpl_137 = (~ and_tmp_7) | mem_inst_request_xbar_xbar_for_3_if_1_mux_28_tmp;
  assign mem_inst_banks_bank_array_impl_data0_rsci_data_in_d = MUX_v_8_8_2(while_req_reg_data_0_lpi_1_dfm_1_mx0,
      while_req_reg_data_1_lpi_1_dfm_1_mx0, while_req_reg_data_2_lpi_1_dfm_1_mx0,
      while_req_reg_data_3_lpi_1_dfm_1_mx0, while_req_reg_data_4_lpi_1_dfm_1_mx0,
      while_req_reg_data_5_lpi_1_dfm_1_mx0, while_req_reg_data_6_lpi_1_dfm_1_mx0,
      while_req_reg_data_7_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_1_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_1_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_1_sva_1});
  assign mem_inst_banks_bank_array_impl_data0_rsci_addr_d = MUX_v_5_8_2(while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_1_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_1_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_1_sva_1});
  assign mem_inst_banks_bank_array_impl_data0_rsci_re_d = ~(and_tmp & and_685_cse
      & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_tmp));
  assign mem_inst_banks_bank_array_impl_data0_rsci_we_d = ~(and_tmp & and_685_cse
      & mem_inst_request_xbar_xbar_for_3_if_1_mux_tmp);
  assign mem_inst_banks_bank_array_impl_data1_rsci_data_in_d = MUX_v_8_8_2(while_req_reg_data_0_lpi_1_dfm_1_mx0,
      while_req_reg_data_1_lpi_1_dfm_1_mx0, while_req_reg_data_2_lpi_1_dfm_1_mx0,
      while_req_reg_data_3_lpi_1_dfm_1_mx0, while_req_reg_data_4_lpi_1_dfm_1_mx0,
      while_req_reg_data_5_lpi_1_dfm_1_mx0, while_req_reg_data_6_lpi_1_dfm_1_mx0,
      while_req_reg_data_7_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_2_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_2_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_2_sva_1});
  assign mem_inst_banks_bank_array_impl_data1_rsci_addr_d = MUX_v_5_8_2(while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_2_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_2_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_2_sva_1});
  assign mem_inst_banks_bank_array_impl_data1_rsci_re_d = ~(and_tmp_1 & and_685_cse
      & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp));
  assign mem_inst_banks_bank_array_impl_data1_rsci_we_d = ~(and_tmp_1 & and_685_cse
      & mem_inst_request_xbar_xbar_for_3_if_1_mux_4_tmp);
  assign mem_inst_banks_bank_array_impl_data2_rsci_data_in_d = MUX_v_8_8_2(while_req_reg_data_0_lpi_1_dfm_1_mx0,
      while_req_reg_data_1_lpi_1_dfm_1_mx0, while_req_reg_data_2_lpi_1_dfm_1_mx0,
      while_req_reg_data_3_lpi_1_dfm_1_mx0, while_req_reg_data_4_lpi_1_dfm_1_mx0,
      while_req_reg_data_5_lpi_1_dfm_1_mx0, while_req_reg_data_6_lpi_1_dfm_1_mx0,
      while_req_reg_data_7_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_3_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_3_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_3_sva_1});
  assign mem_inst_banks_bank_array_impl_data2_rsci_addr_d = MUX_v_5_8_2(while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_3_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_3_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_3_sva_1});
  assign mem_inst_banks_bank_array_impl_data2_rsci_re_d = ~(and_tmp_2 & and_685_cse
      & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp));
  assign mem_inst_banks_bank_array_impl_data2_rsci_we_d = ~(and_tmp_2 & and_685_cse
      & mem_inst_request_xbar_xbar_for_3_if_1_mux_8_tmp);
  assign mem_inst_banks_bank_array_impl_data3_rsci_data_in_d = MUX_v_8_8_2(while_req_reg_data_0_lpi_1_dfm_1_mx0,
      while_req_reg_data_1_lpi_1_dfm_1_mx0, while_req_reg_data_2_lpi_1_dfm_1_mx0,
      while_req_reg_data_3_lpi_1_dfm_1_mx0, while_req_reg_data_4_lpi_1_dfm_1_mx0,
      while_req_reg_data_5_lpi_1_dfm_1_mx0, while_req_reg_data_6_lpi_1_dfm_1_mx0,
      while_req_reg_data_7_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_4_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_4_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_4_sva_1});
  assign mem_inst_banks_bank_array_impl_data3_rsci_addr_d = MUX_v_5_8_2(while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_4_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_4_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_4_sva_1});
  assign mem_inst_banks_bank_array_impl_data3_rsci_re_d = ~(and_tmp_3 & and_685_cse
      & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp));
  assign mem_inst_banks_bank_array_impl_data3_rsci_we_d = ~(and_tmp_3 & and_685_cse
      & mem_inst_request_xbar_xbar_for_3_if_1_mux_12_tmp);
  assign mem_inst_banks_bank_array_impl_data4_rsci_data_in_d = MUX_v_8_8_2(while_req_reg_data_0_lpi_1_dfm_1_mx0,
      while_req_reg_data_1_lpi_1_dfm_1_mx0, while_req_reg_data_2_lpi_1_dfm_1_mx0,
      while_req_reg_data_3_lpi_1_dfm_1_mx0, while_req_reg_data_4_lpi_1_dfm_1_mx0,
      while_req_reg_data_5_lpi_1_dfm_1_mx0, while_req_reg_data_6_lpi_1_dfm_1_mx0,
      while_req_reg_data_7_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_5_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_5_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_5_sva_1});
  assign mem_inst_banks_bank_array_impl_data4_rsci_addr_d = MUX_v_5_8_2(while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_5_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_5_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_5_sva_1});
  assign mem_inst_banks_bank_array_impl_data4_rsci_re_d = ~(and_tmp_4 & and_685_cse
      & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp));
  assign mem_inst_banks_bank_array_impl_data4_rsci_we_d = ~(and_tmp_4 & and_685_cse
      & mem_inst_request_xbar_xbar_for_3_if_1_mux_16_tmp);
  assign mem_inst_banks_bank_array_impl_data5_rsci_data_in_d = MUX_v_8_8_2(while_req_reg_data_0_lpi_1_dfm_1_mx0,
      while_req_reg_data_1_lpi_1_dfm_1_mx0, while_req_reg_data_2_lpi_1_dfm_1_mx0,
      while_req_reg_data_3_lpi_1_dfm_1_mx0, while_req_reg_data_4_lpi_1_dfm_1_mx0,
      while_req_reg_data_5_lpi_1_dfm_1_mx0, while_req_reg_data_6_lpi_1_dfm_1_mx0,
      while_req_reg_data_7_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_6_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_6_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_6_sva_1});
  assign mem_inst_banks_bank_array_impl_data5_rsci_addr_d = MUX_v_5_8_2(while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_6_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_6_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_6_sva_1});
  assign mem_inst_banks_bank_array_impl_data5_rsci_re_d = ~(and_tmp_5 & and_685_cse
      & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp));
  assign mem_inst_banks_bank_array_impl_data5_rsci_we_d = ~(and_tmp_5 & and_685_cse
      & mem_inst_request_xbar_xbar_for_3_if_1_mux_20_tmp);
  assign mem_inst_banks_bank_array_impl_data6_rsci_data_in_d = MUX_v_8_8_2(while_req_reg_data_0_lpi_1_dfm_1_mx0,
      while_req_reg_data_1_lpi_1_dfm_1_mx0, while_req_reg_data_2_lpi_1_dfm_1_mx0,
      while_req_reg_data_3_lpi_1_dfm_1_mx0, while_req_reg_data_4_lpi_1_dfm_1_mx0,
      while_req_reg_data_5_lpi_1_dfm_1_mx0, while_req_reg_data_6_lpi_1_dfm_1_mx0,
      while_req_reg_data_7_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_7_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_7_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_7_sva_1});
  assign mem_inst_banks_bank_array_impl_data6_rsci_addr_d = MUX_v_5_8_2(while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_7_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_7_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_7_sva_1});
  assign mem_inst_banks_bank_array_impl_data6_rsci_re_d = ~(and_tmp_6 & and_685_cse
      & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp));
  assign mem_inst_banks_bank_array_impl_data6_rsci_we_d = ~(and_tmp_6 & and_685_cse
      & mem_inst_request_xbar_xbar_for_3_if_1_mux_24_tmp);
  assign mem_inst_banks_bank_array_impl_data7_rsci_data_in_d = MUX_v_8_8_2(while_req_reg_data_0_lpi_1_dfm_1_mx0,
      while_req_reg_data_1_lpi_1_dfm_1_mx0, while_req_reg_data_2_lpi_1_dfm_1_mx0,
      while_req_reg_data_3_lpi_1_dfm_1_mx0, while_req_reg_data_4_lpi_1_dfm_1_mx0,
      while_req_reg_data_5_lpi_1_dfm_1_mx0, while_req_reg_data_6_lpi_1_dfm_1_mx0,
      while_req_reg_data_7_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_sva_1});
  assign mem_inst_banks_bank_array_impl_data7_rsci_addr_d = MUX_v_5_8_2(while_req_reg_addr_0_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_1_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_2_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_3_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_4_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_5_7_3_lpi_1_dfm_1_mx0, while_req_reg_addr_6_7_3_lpi_1_dfm_1_mx0,
      while_req_reg_addr_7_7_3_lpi_1_dfm_1_mx0, {one_hot_to_bin_8U_3U_for_3_for_1_8_operator_1_false_11_or_psp_sva_1
      , one_hot_to_bin_8U_3U_for_2_for_1_8_operator_1_false_11_or_psp_sva_1 , one_hot_to_bin_8U_3U_for_1_for_1_8_operator_1_false_11_or_psp_sva_1});
  assign mem_inst_banks_bank_array_impl_data7_rsci_re_d = ~(and_tmp_7 & and_685_cse
      & (~ mem_inst_request_xbar_xbar_for_3_if_1_mux_28_tmp));
  assign mem_inst_banks_bank_array_impl_data7_rsci_we_d = ~(and_tmp_7 & and_685_cse
      & mem_inst_request_xbar_xbar_for_3_if_1_mux_28_tmp);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_1_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_1_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0);
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6 & operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5 & operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4 & operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3 & operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2 & operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1 & operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_1_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_1_sva_1);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_1 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_2_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_1 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_1
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_1 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_1 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_1
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_1 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_1 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_1
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_1 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_2_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_1 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_1
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_1 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_1
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_1 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_1
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_1 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_1
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0);
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_1 & operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_1 & operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_1 & operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_1 & operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_1 & operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_1 & operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_1 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_2_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_1 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_1 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_1 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_1 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_1 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_1 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_2_sva_1);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_2 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_3_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_2 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_2
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_2 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_2 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_2
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_2 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_2 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_2
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_2 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_3_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_3_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_2 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_2
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_2 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_2
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_2 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_2
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_2 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_2
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0);
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_14
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_2 & operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_13
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_2 & operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_12
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_2 & operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_11
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_2 & operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_10
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_2 & operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_9
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_2 & operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1;
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_2 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_3_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_6
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_2 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_5
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_2 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_4
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_2 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_3
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_2 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_2
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_2 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1);
  assign mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_1
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_2 & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_3_sva_1);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_3 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_4_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_3 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_3
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_3 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_3 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_3
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_3 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_3 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_3
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_3 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_4_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_4_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_3 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_3
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_3 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_3
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_3 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_3
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_3 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_3
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0);
  assign mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_3 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_4_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_4_sva_1);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_4 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_5_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_4 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_4
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_4 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_4 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_4
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_4 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_4 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_4
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_4 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_5_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_5_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_4 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_4
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_4 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_4
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_4 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_4
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_4 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_4
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0);
  assign mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_4 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_5_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_5_sva_1);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_5 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_6_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_5 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_5
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_5 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_5 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_5
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_5 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_5 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_5
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_5 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_6_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_6_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_5 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_5
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_5 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_5
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_5 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_5
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_5 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_5
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0);
  assign mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_5 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_6_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_6_sva_1);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_6 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_7_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_6 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_6
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_6 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_6 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_6
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_6 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_6 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_6
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_6 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_7_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_7_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_6 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_6
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_6 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_6
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_6 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_6
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_6 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_6
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0);
  assign mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_6 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_7_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_7_sva_1);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_7 = (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_lpi_1_dfm_mx0)
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_6_7 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_7
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_7 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_lpi_1_dfm_mx0
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_5_7 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_7
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_7 = ~(nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_lpi_1_dfm_mx0
      | nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_4_7 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_7
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_7 = nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_0_lpi_1_dfm_mx0
      & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_1_lpi_1_dfm_mx0;
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_3_7 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_7
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_2_7 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_2_7
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_1_7 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_1_7
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0);
  assign Arbiter_8U_Roundrobin_pick_if_1_and_stg_2_0_7 = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_0_7
      & (~ nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0);
  assign mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_wrs_Arbiter_8U_Roundrobin_pick_unrolled_choice_Arbiter_8U_Roundrobin_pick_first_one_idx_1_0_tmp_7
      = Arbiter_8U_Roundrobin_pick_if_1_and_stg_1_3_7 & nvhls_leading_ones_15U_Arbiter_8U_Roundrobin_UnrolledMask_nvhls_nvhls_t_4U_nvuint_t_idx_2_lpi_1_dfm_mx0
      & (~ operator_7_false_operator_7_false_operator_7_false_or_mdf_sva_1);
  assign crossbar_InputSetup_InputType_8U_8U_for_and_20_cse = while_lor_lpi_1_dfm_2
      & (fsm_output[1]);
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      reg_mem_inst_banks_bank_array_impl_data7_rsc_cgo_cse <= 1'b0;
      reg_mem_inst_banks_bank_array_impl_data6_rsc_cgo_cse <= 1'b0;
      reg_mem_inst_banks_bank_array_impl_data5_rsc_cgo_cse <= 1'b0;
      reg_mem_inst_banks_bank_array_impl_data4_rsc_cgo_cse <= 1'b0;
      reg_mem_inst_banks_bank_array_impl_data3_rsc_cgo_cse <= 1'b0;
      reg_mem_inst_banks_bank_array_impl_data2_rsc_cgo_cse <= 1'b0;
      reg_mem_inst_banks_bank_array_impl_data1_rsc_cgo_cse <= 1'b0;
      reg_mem_inst_banks_bank_array_impl_data0_rsc_cgo_cse <= 1'b0;
      reg_rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse <= 1'b0;
      reg_write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse <= 1'b0;
      reg_req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse <= 1'b0;
      while_stage_0_3 <= 1'b0;
      while_stage_0_4 <= 1'b0;
      while_stage_0_5 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_1_1 <= 3'b000;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_1_1 <= 3'b000;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_1_1 <= 3'b000;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_1_1 <= 3'b000;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_1_1 <= 3'b000;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_1_1 <= 3'b000;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_1_1 <= 3'b000;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_1_1 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp ) begin
      reg_mem_inst_banks_bank_array_impl_data7_rsc_cgo_cse <= and_511_rmff;
      reg_mem_inst_banks_bank_array_impl_data6_rsc_cgo_cse <= and_513_rmff;
      reg_mem_inst_banks_bank_array_impl_data5_rsc_cgo_cse <= and_515_rmff;
      reg_mem_inst_banks_bank_array_impl_data4_rsc_cgo_cse <= and_517_rmff;
      reg_mem_inst_banks_bank_array_impl_data3_rsc_cgo_cse <= and_519_rmff;
      reg_mem_inst_banks_bank_array_impl_data2_rsc_cgo_cse <= and_521_rmff;
      reg_mem_inst_banks_bank_array_impl_data1_rsc_cgo_cse <= and_523_rmff;
      reg_mem_inst_banks_bank_array_impl_data0_rsc_cgo_cse <= and_525_rmff;
      reg_rsp_inter_Push_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse <= and_dcpl;
      reg_write_req_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse <= and_231_rmff;
      reg_req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse <= fsm_output[1];
      while_stage_0_3 <= reg_req_inter_PopNB_mioi_ccs_ccore_start_rsc_dat_MemoryRun_psct_cse;
      while_stage_0_4 <= while_stage_0_3;
      while_stage_0_5 <= while_stage_0_4;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_1_1 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_1_1 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_1_1 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_1_1 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_1_1 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_1_1 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_1_1 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_1_1 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp & or_dcpl_1 & and_dcpl_1 & crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1
        ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1_dfm_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1_dfm_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1_dfm_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1_dfm_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1_dfm_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1_dfm_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( crossbar_InputSetup_InputType_8U_8U_for_aelse_and_8_cse ) begin
      crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp & or_dcpl_1 & and_dcpl_1 & crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1
        ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp & or_dcpl_1 & and_dcpl_1 & crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1
        ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp & or_dcpl_1 & and_dcpl_1 & crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1
        ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp & or_dcpl_1 & and_dcpl_1 & crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1
        ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp & or_dcpl_1 & and_dcpl_1 & crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1
        ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp & or_dcpl_1 & and_dcpl_1 & crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1
        ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= 3'b000;
    end
    else if ( rsp_inter_Push_mioi_wen_comp & or_dcpl_1 & and_dcpl_1 & crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1
        ) begin
      crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_2 <= crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_1_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= 8'b00000000;
      mem_inst_load_store_data_out_0_lpi_1_dfm_1 <= 8'b00000000;
      crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= 8'b00000000;
      crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= 8'b00000000;
      crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= 8'b00000000;
      crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= 8'b00000000;
      crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= 8'b00000000;
      crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= 8'b00000000;
    end
    else if ( crossbar_InputSetup_InputType_8U_8U_for_and_7_cse ) begin
      crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
          crossbar_InputSetup_InputType_8U_8U_for_8_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
          or_dcpl_11);
      mem_inst_load_store_data_out_0_lpi_1_dfm_1 <= MUX_v_8_2_2(mem_inst_load_store_data_out_0_lpi_1_dfm_2,
          mem_inst_load_store_data_out_0_lpi_1_dfm_1, or_dcpl_11);
      crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
          crossbar_InputSetup_InputType_8U_8U_for_7_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
          or_dcpl_11);
      crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
          crossbar_InputSetup_InputType_8U_8U_for_2_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
          or_dcpl_11);
      crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
          crossbar_InputSetup_InputType_8U_8U_for_6_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
          or_dcpl_11);
      crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
          crossbar_InputSetup_InputType_8U_8U_for_3_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
          or_dcpl_11);
      crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
          crossbar_InputSetup_InputType_8U_8U_for_5_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
          or_dcpl_11);
      crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1
          <= MUX_v_8_2_2(crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_2,
          crossbar_InputSetup_InputType_8U_8U_for_4_slc_mem_inst_load_store_data_in_8_7_0_pmx_lpi_1_dfm_1,
          or_dcpl_11);
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1_dfm_1_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1_dfm_1_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1_dfm_1_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1_dfm_1_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1_dfm_1_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1_dfm_1_2 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1_dfm_1_2 <= 1'b0;
    end
    else if ( crossbar_InputSetup_InputType_8U_8U_for_aelse_and_16_cse ) begin
      crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1_dfm_1_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1_dfm_1_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1_dfm_1_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1_dfm_1_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1_dfm_1_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1_dfm_1_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1;
      crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1_dfm_1_2 <= crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_asn_mdf_sva_st_1_3 <= 1'b0;
      while_lor_lpi_1_dfm_2 <= 1'b0;
    end
    else if ( while_and_itm ) begin
      while_asn_mdf_sva_st_1_3 <= while_asn_mdf_sva_st_1_2;
      while_lor_lpi_1_dfm_2 <= while_lor_lpi_1_dfm_st_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= 1'b0;
      mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= 1'b0;
      mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= 1'b0;
      mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= 1'b0;
      mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= 1'b0;
      mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= 1'b0;
      mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= 1'b0;
      mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= 1'b0;
    end
    else if ( mem_inst_request_xbar_xbar_for_3_and_cse ) begin
      mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= mem_inst_request_xbar_xbar_for_3_8_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
      mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= mem_inst_request_xbar_xbar_for_3_7_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
      mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= mem_inst_request_xbar_xbar_for_3_6_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
      mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= mem_inst_request_xbar_xbar_for_3_5_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
      mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= mem_inst_request_xbar_xbar_for_3_4_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
      mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= mem_inst_request_xbar_xbar_for_3_3_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
      mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= mem_inst_request_xbar_xbar_for_3_2_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
      mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_st_1_1
          <= mem_inst_request_xbar_xbar_for_3_1_mem_inst_request_xbar_xbar_for_3_if_1_operator_8_false_1_or_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_lor_lpi_1_dfm_st_1 <= 1'b0;
      while_asn_mdf_sva_st_1_2 <= 1'b0;
    end
    else if ( while_oelse_and_1_cse ) begin
      while_lor_lpi_1_dfm_st_1 <= while_if_1_while_if_1_or_tmp;
      while_asn_mdf_sva_st_1_2 <= while_asn_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      while_req_reg_addr_sva_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      while_req_reg_data_sva_1 <= 64'b0000000000000000000000000000000000000000000000000000000000000000;
      while_asn_mdf_sva_1 <= 1'b0;
      while_req_reg_type_val_sva_1 <= 1'b0;
      while_req_reg_valids_sva_1 <= 8'b00000000;
    end
    else if ( while_req_reg_addr_and_cse ) begin
      while_req_reg_addr_sva_1 <= req_inter_PopNB_mioi_data_addr_rsc_z_mxwt;
      while_req_reg_data_sva_1 <= req_inter_PopNB_mioi_data_data_rsc_z_mxwt;
      while_asn_mdf_sva_1 <= req_inter_PopNB_mioi_return_rsc_z_mxwt;
      while_req_reg_type_val_sva_1 <= req_inter_PopNB_mioi_data_type_val_rsc_z_mxwt;
      while_req_reg_valids_sva_1 <= req_inter_PopNB_mioi_data_valids_rsc_z_mxwt;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_arbiters_next_0_1_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_0_3_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_0_4_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_0_2_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_0_5_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_0_6_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_0_7_sva <= 1'b1;
    end
    else if ( mem_inst_request_xbar_arbiters_next_and_cse ) begin
      mem_inst_request_xbar_arbiters_next_0_1_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
          | (~ mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_0_3_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_0_4_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_0_2_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_0_5_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_1_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_0_6_sva <= mem_inst_request_xbar_xbar_for_3_1_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
          | (~ mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_0_7_sva <= ~ mem_inst_request_xbar_xbar_for_3_1_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_arbiters_next_1_1_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_1_3_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_1_4_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_1_2_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_1_5_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_1_6_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_1_7_sva <= 1'b1;
    end
    else if ( mem_inst_request_xbar_arbiters_next_and_7_cse ) begin
      mem_inst_request_xbar_arbiters_next_1_1_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
          | (~ mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_1_3_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_1_4_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_1_2_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_1_5_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_2_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_1_6_sva <= mem_inst_request_xbar_xbar_for_3_2_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
          | (~ mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_1_7_sva <= ~ mem_inst_request_xbar_xbar_for_3_2_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_arbiters_next_2_1_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_2_3_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_2_4_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_2_2_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_2_5_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_2_6_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_2_7_sva <= 1'b1;
    end
    else if ( mem_inst_request_xbar_arbiters_next_and_14_cse ) begin
      mem_inst_request_xbar_arbiters_next_2_1_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
          | (~ mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_2_3_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_2_4_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_2_2_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_2_5_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_3_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_2_6_sva <= mem_inst_request_xbar_xbar_for_3_3_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
          | (~ mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_2_7_sva <= ~ mem_inst_request_xbar_xbar_for_3_3_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_arbiters_next_3_1_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_3_3_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_3_4_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_3_2_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_3_5_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_3_6_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_3_7_sva <= 1'b1;
    end
    else if ( mem_inst_request_xbar_arbiters_next_and_21_cse ) begin
      mem_inst_request_xbar_arbiters_next_3_1_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
          | (~ mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_3_3_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_3_4_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_3_2_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_3_5_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_4_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_3_6_sva <= mem_inst_request_xbar_xbar_for_3_4_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
          | (~ mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_3_7_sva <= ~ mem_inst_request_xbar_xbar_for_3_4_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_arbiters_next_4_1_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_4_3_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_4_4_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_4_2_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_4_5_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_4_6_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_4_7_sva <= 1'b1;
    end
    else if ( mem_inst_request_xbar_arbiters_next_and_28_cse ) begin
      mem_inst_request_xbar_arbiters_next_4_1_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
          | (~ mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_4_3_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_4_4_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_4_2_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_4_5_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_5_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_4_6_sva <= mem_inst_request_xbar_xbar_for_3_5_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
          | (~ mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_4_7_sva <= ~ mem_inst_request_xbar_xbar_for_3_5_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_arbiters_next_5_1_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_5_3_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_5_4_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_5_2_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_5_5_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_5_6_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_5_7_sva <= 1'b1;
    end
    else if ( mem_inst_request_xbar_arbiters_next_and_35_cse ) begin
      mem_inst_request_xbar_arbiters_next_5_1_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
          | (~ mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_5_3_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_5_4_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_5_2_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_5_5_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_6_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_5_6_sva <= mem_inst_request_xbar_xbar_for_3_6_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
          | (~ mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_5_7_sva <= ~ mem_inst_request_xbar_xbar_for_3_6_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_arbiters_next_6_1_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_6_3_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_6_4_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_6_2_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_6_5_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_6_6_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_6_7_sva <= 1'b1;
    end
    else if ( mem_inst_request_xbar_arbiters_next_and_42_cse ) begin
      mem_inst_request_xbar_arbiters_next_6_1_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
          | (~ mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_6_3_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_6_4_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_6_2_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_6_5_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_7_sva_1
          | (~ mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_6_6_sva <= mem_inst_request_xbar_xbar_for_3_7_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
          | (~ mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1);
      mem_inst_request_xbar_arbiters_next_6_7_sva <= ~ mem_inst_request_xbar_xbar_for_3_7_operator_4_false_1_operator_4_false_1_nand_mdf_sva_1;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_request_xbar_arbiters_next_7_1_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_7_3_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_7_4_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_7_2_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_7_5_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_7_6_sva <= 1'b1;
      mem_inst_request_xbar_arbiters_next_7_7_sva <= 1'b1;
    end
    else if ( operator_15_false_and_cse ) begin
      mem_inst_request_xbar_arbiters_next_7_1_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_1
          | Arbiter_8U_Roundrobin_pick_if_1_not_64;
      mem_inst_request_xbar_arbiters_next_7_3_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_4_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_if_1_not_64;
      mem_inst_request_xbar_arbiters_next_7_4_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_3_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_if_1_not_64;
      mem_inst_request_xbar_arbiters_next_7_2_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_5_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_if_1_not_64;
      mem_inst_request_xbar_arbiters_next_7_5_sva <= Arbiter_8U_Roundrobin_pick_if_1_if_for_2_Arbiter_8U_Roundrobin_pick_if_1_if_for_or_1_cse_sva_1
          | Arbiter_8U_Roundrobin_pick_if_1_not_64;
      mem_inst_request_xbar_arbiters_next_7_6_sva <= mem_inst_request_xbar_xbar_for_3_8_Arbiter_8U_Roundrobin_pick_if_1_temp2_or_tmp_6
          | Arbiter_8U_Roundrobin_pick_if_1_not_64;
      mem_inst_request_xbar_arbiters_next_7_7_sva <= Arbiter_8U_Roundrobin_pick_if_1_not_64;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1 <= 1'b0;
      crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1 <= 1'b0;
    end
    else if ( crossbar_InputSetup_InputType_8U_8U_for_aelse_and_cse ) begin
      crossbar_InputSetup_InputType_8U_8U_for_land_7_lpi_1 <= (crossbar_InputSetup_InputType_8U_8U_for_mux_27_nl)
          & mem_inst_load_store_valid_src_6_lpi_1_dfm_7_mx0;
      crossbar_InputSetup_InputType_8U_8U_for_land_6_lpi_1 <= (crossbar_InputSetup_InputType_8U_8U_for_mux_25_nl)
          & mem_inst_load_store_valid_src_5_lpi_1_dfm_7_mx0;
      crossbar_InputSetup_InputType_8U_8U_for_land_5_lpi_1 <= (crossbar_InputSetup_InputType_8U_8U_for_mux_23_nl)
          & mem_inst_load_store_valid_src_4_lpi_1_dfm_7_mx0;
      crossbar_InputSetup_InputType_8U_8U_for_land_4_lpi_1 <= (crossbar_InputSetup_InputType_8U_8U_for_mux_21_nl)
          & mem_inst_load_store_valid_src_3_lpi_1_dfm_7_mx0;
      crossbar_InputSetup_InputType_8U_8U_for_land_3_lpi_1 <= (crossbar_InputSetup_InputType_8U_8U_for_mux_19_nl)
          & mem_inst_load_store_valid_src_2_lpi_1_dfm_7_mx0;
      crossbar_InputSetup_InputType_8U_8U_for_land_2_lpi_1 <= (crossbar_InputSetup_InputType_8U_8U_for_mux_17_nl)
          & mem_inst_load_store_valid_src_1_lpi_1_dfm_7_mx0;
      crossbar_InputSetup_InputType_8U_8U_for_land_1_lpi_1 <= (crossbar_InputSetup_InputType_8U_8U_for_mux_14_nl)
          & mem_inst_load_store_valid_src_0_lpi_1_dfm_7_mx0;
      crossbar_InputSetup_InputType_8U_8U_for_land_lpi_1_dfm_1 <= (crossbar_InputSetup_InputType_8U_8U_for_mux_29_nl)
          & mem_inst_load_store_valid_src_7_lpi_1_dfm_7_mx0;
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_1_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_1_1_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_2_1_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_3_1_sva <= 1'b0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_ftd <=
          1'b0;
    end
    else if ( mem_inst_load_store_for_4_if_and_104_cse ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_1_sva <= mem_inst_load_store_for_4_if_and_stg_1_0_1_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_1_1_sva <= mem_inst_load_store_for_4_if_and_stg_1_1_1_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_2_1_sva <= mem_inst_load_store_for_4_if_and_stg_1_2_1_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_3_1_sva <= mem_inst_load_store_for_4_if_and_stg_1_3_1_sva_mx0w0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_ftd <=
          mem_inst_request_xbar_run_1_output_data_input_chan_1_lpi_1_dfm_1_mx0w0[2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_2_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_1_2_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_2_2_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_3_2_sva <= 1'b0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_ftd <=
          1'b0;
    end
    else if ( mem_inst_load_store_for_4_if_and_108_cse ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_2_sva <= mem_inst_load_store_for_4_if_and_stg_1_0_2_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_1_2_sva <= mem_inst_load_store_for_4_if_and_stg_1_1_2_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_2_2_sva <= mem_inst_load_store_for_4_if_and_stg_1_2_2_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_3_2_sva <= mem_inst_load_store_for_4_if_and_stg_1_3_2_sva_mx0w0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_ftd <=
          mem_inst_request_xbar_run_1_output_data_input_chan_2_lpi_1_dfm_1_mx0w0[2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_3_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_1_3_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_2_3_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_3_3_sva <= 1'b0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_ftd <=
          1'b0;
    end
    else if ( mem_inst_load_store_for_4_if_and_112_cse ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_3_sva <= mem_inst_load_store_for_4_if_and_stg_1_0_3_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_1_3_sva <= mem_inst_load_store_for_4_if_and_stg_1_1_3_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_2_3_sva <= mem_inst_load_store_for_4_if_and_stg_1_2_3_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_3_3_sva <= mem_inst_load_store_for_4_if_and_stg_1_3_3_sva_mx0w0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_ftd <=
          mem_inst_request_xbar_run_1_output_data_input_chan_3_lpi_1_dfm_1_mx0w0[2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_4_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_1_4_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_2_4_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_3_4_sva <= 1'b0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_ftd <=
          1'b0;
    end
    else if ( mem_inst_load_store_for_4_if_and_116_cse ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_4_sva <= mem_inst_load_store_for_4_if_and_stg_1_0_4_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_1_4_sva <= mem_inst_load_store_for_4_if_and_stg_1_1_4_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_2_4_sva <= mem_inst_load_store_for_4_if_and_stg_1_2_4_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_3_4_sva <= mem_inst_load_store_for_4_if_and_stg_1_3_4_sva_mx0w0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_ftd <=
          mem_inst_request_xbar_run_1_output_data_input_chan_4_lpi_1_dfm_1_mx0w0[2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_5_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_1_5_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_2_5_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_3_5_sva <= 1'b0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_ftd <=
          1'b0;
    end
    else if ( mem_inst_load_store_for_4_if_and_120_cse ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_5_sva <= mem_inst_load_store_for_4_if_and_stg_1_0_5_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_1_5_sva <= mem_inst_load_store_for_4_if_and_stg_1_1_5_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_2_5_sva <= mem_inst_load_store_for_4_if_and_stg_1_2_5_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_3_5_sva <= mem_inst_load_store_for_4_if_and_stg_1_3_5_sva_mx0w0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_ftd <=
          mem_inst_request_xbar_run_1_output_data_input_chan_5_lpi_1_dfm_1_mx0w0[2];
    end
  end
  always @(posedge clk or negedge rst) begin
    if ( ~ rst ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_6_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_1_6_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_2_6_sva <= 1'b0;
      mem_inst_load_store_for_4_if_and_stg_1_3_6_sva <= 1'b0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_ftd <=
          1'b0;
    end
    else if ( mem_inst_load_store_for_4_if_and_124_cse ) begin
      mem_inst_load_store_for_4_if_and_stg_1_0_6_sva <= mem_inst_load_store_for_4_if_and_stg_1_0_6_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_1_6_sva <= mem_inst_load_store_for_4_if_and_stg_1_1_6_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_2_6_sva <= mem_inst_load_store_for_4_if_and_stg_1_2_6_sva_mx0w0;
      mem_inst_load_store_for_4_if_and_stg_1_3_6_sva <= mem_inst_load_store_for_4_if_and_stg_1_3_6_sva_mx0w0;
      reg_mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_ftd <=
          mem_inst_request_xbar_run_1_output_data_input_chan_6_lpi_1_dfm_1_mx0w0[2];
    end
  end
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_27_nl = MUX_s_1_8_2(mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1, crossbar_InputSetup_InputType_8U_8U_source_tmp_7_lpi_1_dfm_1);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_25_nl = MUX_s_1_8_2(mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1, crossbar_InputSetup_InputType_8U_8U_source_tmp_6_lpi_1_dfm_1);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_23_nl = MUX_s_1_8_2(mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1, crossbar_InputSetup_InputType_8U_8U_source_tmp_5_lpi_1_dfm_1);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_21_nl = MUX_s_1_8_2(mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1, crossbar_InputSetup_InputType_8U_8U_source_tmp_4_lpi_1_dfm_1);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_19_nl = MUX_s_1_8_2(mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1, crossbar_InputSetup_InputType_8U_8U_source_tmp_3_lpi_1_dfm_1);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_17_nl = MUX_s_1_8_2(mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1, crossbar_InputSetup_InputType_8U_8U_source_tmp_2_lpi_1_dfm_1);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_14_nl = MUX_s_1_8_2(mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1, crossbar_InputSetup_InputType_8U_8U_source_tmp_1_lpi_1_dfm_1);
  assign crossbar_InputSetup_InputType_8U_8U_for_mux_29_nl = MUX_s_1_8_2(mem_inst_load_store_bank_rsp_valid_0_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_1_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_2_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_3_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_4_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_5_lpi_1_dfm_1, mem_inst_load_store_bank_rsp_valid_6_lpi_1_dfm_1,
      mem_inst_load_store_bank_rsp_valid_7_lpi_1_dfm_1, crossbar_InputSetup_InputType_8U_8U_source_tmp_lpi_1_dfm_1);

  function automatic [0:0] MUX1HOT_s_1_1_2;
    input [0:0] input_0;
    input [0:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    MUX1HOT_s_1_1_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_4_2;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [3:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    MUX1HOT_s_1_4_2 = result;
  end
  endfunction


  function automatic [0:0] MUX1HOT_s_1_7_2;
    input [0:0] input_6;
    input [0:0] input_5;
    input [0:0] input_4;
    input [0:0] input_3;
    input [0:0] input_2;
    input [0:0] input_1;
    input [0:0] input_0;
    input [6:0] sel;
    reg [0:0] result;
  begin
    result = input_0 & {1{sel[0]}};
    result = result | ( input_1 & {1{sel[1]}});
    result = result | ( input_2 & {1{sel[2]}});
    result = result | ( input_3 & {1{sel[3]}});
    result = result | ( input_4 & {1{sel[4]}});
    result = result | ( input_5 & {1{sel[5]}});
    result = result | ( input_6 & {1{sel[6]}});
    MUX1HOT_s_1_7_2 = result;
  end
  endfunction


  function automatic [2:0] MUX1HOT_v_3_7_2;
    input [2:0] input_6;
    input [2:0] input_5;
    input [2:0] input_4;
    input [2:0] input_3;
    input [2:0] input_2;
    input [2:0] input_1;
    input [2:0] input_0;
    input [6:0] sel;
    reg [2:0] result;
  begin
    result = input_0 & {3{sel[0]}};
    result = result | ( input_1 & {3{sel[1]}});
    result = result | ( input_2 & {3{sel[2]}});
    result = result | ( input_3 & {3{sel[3]}});
    result = result | ( input_4 & {3{sel[4]}});
    result = result | ( input_5 & {3{sel[5]}});
    result = result | ( input_6 & {3{sel[6]}});
    MUX1HOT_v_3_7_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_2_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function automatic [0:0] MUX_s_1_8_2;
    input [0:0] input_0;
    input [0:0] input_1;
    input [0:0] input_2;
    input [0:0] input_3;
    input [0:0] input_4;
    input [0:0] input_5;
    input [0:0] input_6;
    input [0:0] input_7;
    input [2:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_s_1_8_2 = result;
  end
  endfunction


  function automatic [1:0] MUX_v_2_2_2;
    input [1:0] input_0;
    input [1:0] input_1;
    input [0:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_2_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_2_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function automatic [2:0] MUX_v_3_8_2;
    input [2:0] input_0;
    input [2:0] input_1;
    input [2:0] input_2;
    input [2:0] input_3;
    input [2:0] input_4;
    input [2:0] input_5;
    input [2:0] input_6;
    input [2:0] input_7;
    input [2:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_3_8_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_2_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [0:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_5_2_2 = result;
  end
  endfunction


  function automatic [4:0] MUX_v_5_8_2;
    input [4:0] input_0;
    input [4:0] input_1;
    input [4:0] input_2;
    input [4:0] input_3;
    input [4:0] input_4;
    input [4:0] input_5;
    input [4:0] input_6;
    input [4:0] input_7;
    input [2:0] sel;
    reg [4:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_5_8_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_2_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [0:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = input_0;
      end
      default : begin
        result = input_1;
      end
    endcase
    MUX_v_8_2_2 = result;
  end
  endfunction


  function automatic [7:0] MUX_v_8_8_2;
    input [7:0] input_0;
    input [7:0] input_1;
    input [7:0] input_2;
    input [7:0] input_3;
    input [7:0] input_4;
    input [7:0] input_5;
    input [7:0] input_6;
    input [7:0] input_7;
    input [2:0] sel;
    reg [7:0] result;
  begin
    case (sel)
      3'b000 : begin
        result = input_0;
      end
      3'b001 : begin
        result = input_1;
      end
      3'b010 : begin
        result = input_2;
      end
      3'b011 : begin
        result = input_3;
      end
      3'b100 : begin
        result = input_4;
      end
      3'b101 : begin
        result = input_5;
      end
      3'b110 : begin
        result = input_6;
      end
      default : begin
        result = input_7;
      end
    endcase
    MUX_v_8_8_2 = result;
  end
  endfunction


  function automatic [1:0] signext_2_1;
    input [0:0] vector;
  begin
    signext_2_1= {{1{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function automatic [2:0] signext_3_2;
    input [1:0] vector;
  begin
    signext_3_2= {{1{vector[1]}}, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysPE
// ------------------------------------------------------------------


module SysPE (
  clk, rst, weight_in_val, weight_in_rdy, weight_in_msg, act_in_val, act_in_rdy,
      act_in_msg, accum_in_val, accum_in_rdy, accum_in_msg, act_out_val, act_out_rdy,
      act_out_msg, accum_out_val, accum_out_rdy, accum_out_msg, weight_out_val, weight_out_rdy,
      weight_out_msg
);
  input clk;
  input rst;
  input weight_in_val;
  output weight_in_rdy;
  input [7:0] weight_in_msg;
  input act_in_val;
  output act_in_rdy;
  input [7:0] act_in_msg;
  input accum_in_val;
  output accum_in_rdy;
  input [31:0] accum_in_msg;
  output act_out_val;
  input act_out_rdy;
  output [7:0] act_out_msg;
  output accum_out_val;
  input accum_out_rdy;
  output [31:0] accum_out_msg;
  output weight_out_val;
  input weight_out_rdy;
  output [7:0] weight_out_msg;



  // Interconnect Declarations for Component Instantiations 
  SysPE_PERun SysPE_PERun_inst (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_val),
      .weight_in_rdy(weight_in_rdy),
      .weight_in_msg(weight_in_msg),
      .act_in_val(act_in_val),
      .act_in_rdy(act_in_rdy),
      .act_in_msg(act_in_msg),
      .accum_in_val(accum_in_val),
      .accum_in_rdy(accum_in_rdy),
      .accum_in_msg(accum_in_msg),
      .act_out_val(act_out_val),
      .act_out_rdy(act_out_rdy),
      .act_out_msg(act_out_msg),
      .accum_out_val(accum_out_val),
      .accum_out_rdy(accum_out_rdy),
      .accum_out_msg(accum_out_msg),
      .weight_out_val(weight_out_val),
      .weight_out_rdy(weight_out_rdy),
      .weight_out_msg(weight_out_msg)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    InputSetup
// ------------------------------------------------------------------


module InputSetup (
  clk, rst, write_req_val, write_req_rdy, write_req_msg, start_val, start_rdy, start_msg,
      act_in_vec_0_val, act_in_vec_1_val, act_in_vec_2_val, act_in_vec_3_val, act_in_vec_4_val,
      act_in_vec_5_val, act_in_vec_6_val, act_in_vec_7_val, act_in_vec_0_rdy, act_in_vec_1_rdy,
      act_in_vec_2_rdy, act_in_vec_3_rdy, act_in_vec_4_rdy, act_in_vec_5_rdy, act_in_vec_6_rdy,
      act_in_vec_7_rdy, act_in_vec_0_msg, act_in_vec_1_msg, act_in_vec_2_msg, act_in_vec_3_msg,
      act_in_vec_4_msg, act_in_vec_5_msg, act_in_vec_6_msg, act_in_vec_7_msg
);
  input clk;
  input rst;
  input write_req_val;
  output write_req_rdy;
  input [68:0] write_req_msg;
  input start_val;
  output start_rdy;
  input [5:0] start_msg;
  output act_in_vec_0_val;
  output act_in_vec_1_val;
  output act_in_vec_2_val;
  output act_in_vec_3_val;
  output act_in_vec_4_val;
  output act_in_vec_5_val;
  output act_in_vec_6_val;
  output act_in_vec_7_val;
  input act_in_vec_0_rdy;
  input act_in_vec_1_rdy;
  input act_in_vec_2_rdy;
  input act_in_vec_3_rdy;
  input act_in_vec_4_rdy;
  input act_in_vec_5_rdy;
  input act_in_vec_6_rdy;
  input act_in_vec_7_rdy;
  output [7:0] act_in_vec_0_msg;
  output [7:0] act_in_vec_1_msg;
  output [7:0] act_in_vec_2_msg;
  output [7:0] act_in_vec_3_msg;
  output [7:0] act_in_vec_4_msg;
  output [7:0] act_in_vec_5_msg;
  output [7:0] act_in_vec_6_msg;
  output [7:0] act_in_vec_7_msg;


  // Interconnect Declarations
  wire req_inter_val;
  wire req_inter_rdy;
  wire [136:0] req_inter_msg;
  wire rsp_inter_val;
  wire rsp_inter_rdy;
  wire [71:0] rsp_inter_msg;
  wire [7:0] mem_inst_banks_bank_array_impl_data0_rsci_data_in_d;
  wire [4:0] mem_inst_banks_bank_array_impl_data0_rsci_addr_d;
  wire mem_inst_banks_bank_array_impl_data0_rsci_re_d;
  wire mem_inst_banks_bank_array_impl_data0_rsci_we_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data0_rsci_data_out_d;
  wire mem_inst_banks_bank_array_impl_data0_rsci_en_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data1_rsci_data_in_d;
  wire [4:0] mem_inst_banks_bank_array_impl_data1_rsci_addr_d;
  wire mem_inst_banks_bank_array_impl_data1_rsci_re_d;
  wire mem_inst_banks_bank_array_impl_data1_rsci_we_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data1_rsci_data_out_d;
  wire mem_inst_banks_bank_array_impl_data1_rsci_en_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data2_rsci_data_in_d;
  wire [4:0] mem_inst_banks_bank_array_impl_data2_rsci_addr_d;
  wire mem_inst_banks_bank_array_impl_data2_rsci_re_d;
  wire mem_inst_banks_bank_array_impl_data2_rsci_we_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data2_rsci_data_out_d;
  wire mem_inst_banks_bank_array_impl_data2_rsci_en_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data3_rsci_data_in_d;
  wire [4:0] mem_inst_banks_bank_array_impl_data3_rsci_addr_d;
  wire mem_inst_banks_bank_array_impl_data3_rsci_re_d;
  wire mem_inst_banks_bank_array_impl_data3_rsci_we_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data3_rsci_data_out_d;
  wire mem_inst_banks_bank_array_impl_data3_rsci_en_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data4_rsci_data_in_d;
  wire [4:0] mem_inst_banks_bank_array_impl_data4_rsci_addr_d;
  wire mem_inst_banks_bank_array_impl_data4_rsci_re_d;
  wire mem_inst_banks_bank_array_impl_data4_rsci_we_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data4_rsci_data_out_d;
  wire mem_inst_banks_bank_array_impl_data4_rsci_en_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data5_rsci_data_in_d;
  wire [4:0] mem_inst_banks_bank_array_impl_data5_rsci_addr_d;
  wire mem_inst_banks_bank_array_impl_data5_rsci_re_d;
  wire mem_inst_banks_bank_array_impl_data5_rsci_we_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data5_rsci_data_out_d;
  wire mem_inst_banks_bank_array_impl_data5_rsci_en_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data6_rsci_data_in_d;
  wire [4:0] mem_inst_banks_bank_array_impl_data6_rsci_addr_d;
  wire mem_inst_banks_bank_array_impl_data6_rsci_re_d;
  wire mem_inst_banks_bank_array_impl_data6_rsci_we_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data6_rsci_data_out_d;
  wire mem_inst_banks_bank_array_impl_data6_rsci_en_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data7_rsci_data_in_d;
  wire [4:0] mem_inst_banks_bank_array_impl_data7_rsci_addr_d;
  wire mem_inst_banks_bank_array_impl_data7_rsci_re_d;
  wire mem_inst_banks_bank_array_impl_data7_rsci_we_d;
  wire [7:0] mem_inst_banks_bank_array_impl_data7_rsci_data_out_d;
  wire mem_inst_banks_bank_array_impl_data7_rsci_en_d;
  wire mem_inst_banks_bank_array_impl_data0_rsc_en;
  wire [7:0] mem_inst_banks_bank_array_impl_data0_rsc_data_out;
  wire mem_inst_banks_bank_array_impl_data0_rsc_we;
  wire mem_inst_banks_bank_array_impl_data0_rsc_re;
  wire [4:0] mem_inst_banks_bank_array_impl_data0_rsc_addr;
  wire [7:0] mem_inst_banks_bank_array_impl_data0_rsc_data_in;
  wire mem_inst_banks_bank_array_impl_data1_rsc_en;
  wire [7:0] mem_inst_banks_bank_array_impl_data1_rsc_data_out;
  wire mem_inst_banks_bank_array_impl_data1_rsc_we;
  wire mem_inst_banks_bank_array_impl_data1_rsc_re;
  wire [4:0] mem_inst_banks_bank_array_impl_data1_rsc_addr;
  wire [7:0] mem_inst_banks_bank_array_impl_data1_rsc_data_in;
  wire mem_inst_banks_bank_array_impl_data2_rsc_en;
  wire [7:0] mem_inst_banks_bank_array_impl_data2_rsc_data_out;
  wire mem_inst_banks_bank_array_impl_data2_rsc_we;
  wire mem_inst_banks_bank_array_impl_data2_rsc_re;
  wire [4:0] mem_inst_banks_bank_array_impl_data2_rsc_addr;
  wire [7:0] mem_inst_banks_bank_array_impl_data2_rsc_data_in;
  wire mem_inst_banks_bank_array_impl_data3_rsc_en;
  wire [7:0] mem_inst_banks_bank_array_impl_data3_rsc_data_out;
  wire mem_inst_banks_bank_array_impl_data3_rsc_we;
  wire mem_inst_banks_bank_array_impl_data3_rsc_re;
  wire [4:0] mem_inst_banks_bank_array_impl_data3_rsc_addr;
  wire [7:0] mem_inst_banks_bank_array_impl_data3_rsc_data_in;
  wire mem_inst_banks_bank_array_impl_data4_rsc_en;
  wire [7:0] mem_inst_banks_bank_array_impl_data4_rsc_data_out;
  wire mem_inst_banks_bank_array_impl_data4_rsc_we;
  wire mem_inst_banks_bank_array_impl_data4_rsc_re;
  wire [4:0] mem_inst_banks_bank_array_impl_data4_rsc_addr;
  wire [7:0] mem_inst_banks_bank_array_impl_data4_rsc_data_in;
  wire mem_inst_banks_bank_array_impl_data5_rsc_en;
  wire [7:0] mem_inst_banks_bank_array_impl_data5_rsc_data_out;
  wire mem_inst_banks_bank_array_impl_data5_rsc_we;
  wire mem_inst_banks_bank_array_impl_data5_rsc_re;
  wire [4:0] mem_inst_banks_bank_array_impl_data5_rsc_addr;
  wire [7:0] mem_inst_banks_bank_array_impl_data5_rsc_data_in;
  wire mem_inst_banks_bank_array_impl_data6_rsc_en;
  wire [7:0] mem_inst_banks_bank_array_impl_data6_rsc_data_out;
  wire mem_inst_banks_bank_array_impl_data6_rsc_we;
  wire mem_inst_banks_bank_array_impl_data6_rsc_re;
  wire [4:0] mem_inst_banks_bank_array_impl_data6_rsc_addr;
  wire [7:0] mem_inst_banks_bank_array_impl_data6_rsc_data_in;
  wire mem_inst_banks_bank_array_impl_data7_rsc_en;
  wire [7:0] mem_inst_banks_bank_array_impl_data7_rsc_data_out;
  wire mem_inst_banks_bank_array_impl_data7_rsc_we;
  wire mem_inst_banks_bank_array_impl_data7_rsc_re;
  wire [4:0] mem_inst_banks_bank_array_impl_data7_rsc_addr;
  wire [7:0] mem_inst_banks_bank_array_impl_data7_rsc_data_in;


  // Interconnect Declarations for Component Instantiations 
  ram_sync_single_be #(.ram_id(32'sd297),
  .words(32'sd32),
  .width(32'sd8),
  .addr_width(32'sd5),
  .a_reset_active(32'sd0),
  .s_reset_active(32'sd0),
  .enable_active(32'sd0),
  .re_active(32'sd0),
  .we_active(32'sd0),
  .num_byte_enables(32'sd1),
  .clock_edge(32'sd1),
  .no_of_RAM_readwrite_port(32'sd1)) mem_inst_banks_bank_array_impl_data0_rsc_comp
      (
      .data_in(mem_inst_banks_bank_array_impl_data0_rsc_data_in),
      .addr(mem_inst_banks_bank_array_impl_data0_rsc_addr),
      .re(mem_inst_banks_bank_array_impl_data0_rsc_re),
      .we(mem_inst_banks_bank_array_impl_data0_rsc_we),
      .data_out(mem_inst_banks_bank_array_impl_data0_rsc_data_out),
      .clk(clk),
      .a_rst(rst),
      .s_rst(1'b1),
      .en(mem_inst_banks_bank_array_impl_data0_rsc_en)
    );
  ram_sync_single_be #(.ram_id(32'sd298),
  .words(32'sd32),
  .width(32'sd8),
  .addr_width(32'sd5),
  .a_reset_active(32'sd0),
  .s_reset_active(32'sd0),
  .enable_active(32'sd0),
  .re_active(32'sd0),
  .we_active(32'sd0),
  .num_byte_enables(32'sd1),
  .clock_edge(32'sd1),
  .no_of_RAM_readwrite_port(32'sd1)) mem_inst_banks_bank_array_impl_data1_rsc_comp
      (
      .data_in(mem_inst_banks_bank_array_impl_data1_rsc_data_in),
      .addr(mem_inst_banks_bank_array_impl_data1_rsc_addr),
      .re(mem_inst_banks_bank_array_impl_data1_rsc_re),
      .we(mem_inst_banks_bank_array_impl_data1_rsc_we),
      .data_out(mem_inst_banks_bank_array_impl_data1_rsc_data_out),
      .clk(clk),
      .a_rst(rst),
      .s_rst(1'b1),
      .en(mem_inst_banks_bank_array_impl_data1_rsc_en)
    );
  ram_sync_single_be #(.ram_id(32'sd299),
  .words(32'sd32),
  .width(32'sd8),
  .addr_width(32'sd5),
  .a_reset_active(32'sd0),
  .s_reset_active(32'sd0),
  .enable_active(32'sd0),
  .re_active(32'sd0),
  .we_active(32'sd0),
  .num_byte_enables(32'sd1),
  .clock_edge(32'sd1),
  .no_of_RAM_readwrite_port(32'sd1)) mem_inst_banks_bank_array_impl_data2_rsc_comp
      (
      .data_in(mem_inst_banks_bank_array_impl_data2_rsc_data_in),
      .addr(mem_inst_banks_bank_array_impl_data2_rsc_addr),
      .re(mem_inst_banks_bank_array_impl_data2_rsc_re),
      .we(mem_inst_banks_bank_array_impl_data2_rsc_we),
      .data_out(mem_inst_banks_bank_array_impl_data2_rsc_data_out),
      .clk(clk),
      .a_rst(rst),
      .s_rst(1'b1),
      .en(mem_inst_banks_bank_array_impl_data2_rsc_en)
    );
  ram_sync_single_be #(.ram_id(32'sd300),
  .words(32'sd32),
  .width(32'sd8),
  .addr_width(32'sd5),
  .a_reset_active(32'sd0),
  .s_reset_active(32'sd0),
  .enable_active(32'sd0),
  .re_active(32'sd0),
  .we_active(32'sd0),
  .num_byte_enables(32'sd1),
  .clock_edge(32'sd1),
  .no_of_RAM_readwrite_port(32'sd1)) mem_inst_banks_bank_array_impl_data3_rsc_comp
      (
      .data_in(mem_inst_banks_bank_array_impl_data3_rsc_data_in),
      .addr(mem_inst_banks_bank_array_impl_data3_rsc_addr),
      .re(mem_inst_banks_bank_array_impl_data3_rsc_re),
      .we(mem_inst_banks_bank_array_impl_data3_rsc_we),
      .data_out(mem_inst_banks_bank_array_impl_data3_rsc_data_out),
      .clk(clk),
      .a_rst(rst),
      .s_rst(1'b1),
      .en(mem_inst_banks_bank_array_impl_data3_rsc_en)
    );
  ram_sync_single_be #(.ram_id(32'sd301),
  .words(32'sd32),
  .width(32'sd8),
  .addr_width(32'sd5),
  .a_reset_active(32'sd0),
  .s_reset_active(32'sd0),
  .enable_active(32'sd0),
  .re_active(32'sd0),
  .we_active(32'sd0),
  .num_byte_enables(32'sd1),
  .clock_edge(32'sd1),
  .no_of_RAM_readwrite_port(32'sd1)) mem_inst_banks_bank_array_impl_data4_rsc_comp
      (
      .data_in(mem_inst_banks_bank_array_impl_data4_rsc_data_in),
      .addr(mem_inst_banks_bank_array_impl_data4_rsc_addr),
      .re(mem_inst_banks_bank_array_impl_data4_rsc_re),
      .we(mem_inst_banks_bank_array_impl_data4_rsc_we),
      .data_out(mem_inst_banks_bank_array_impl_data4_rsc_data_out),
      .clk(clk),
      .a_rst(rst),
      .s_rst(1'b1),
      .en(mem_inst_banks_bank_array_impl_data4_rsc_en)
    );
  ram_sync_single_be #(.ram_id(32'sd302),
  .words(32'sd32),
  .width(32'sd8),
  .addr_width(32'sd5),
  .a_reset_active(32'sd0),
  .s_reset_active(32'sd0),
  .enable_active(32'sd0),
  .re_active(32'sd0),
  .we_active(32'sd0),
  .num_byte_enables(32'sd1),
  .clock_edge(32'sd1),
  .no_of_RAM_readwrite_port(32'sd1)) mem_inst_banks_bank_array_impl_data5_rsc_comp
      (
      .data_in(mem_inst_banks_bank_array_impl_data5_rsc_data_in),
      .addr(mem_inst_banks_bank_array_impl_data5_rsc_addr),
      .re(mem_inst_banks_bank_array_impl_data5_rsc_re),
      .we(mem_inst_banks_bank_array_impl_data5_rsc_we),
      .data_out(mem_inst_banks_bank_array_impl_data5_rsc_data_out),
      .clk(clk),
      .a_rst(rst),
      .s_rst(1'b1),
      .en(mem_inst_banks_bank_array_impl_data5_rsc_en)
    );
  ram_sync_single_be #(.ram_id(32'sd303),
  .words(32'sd32),
  .width(32'sd8),
  .addr_width(32'sd5),
  .a_reset_active(32'sd0),
  .s_reset_active(32'sd0),
  .enable_active(32'sd0),
  .re_active(32'sd0),
  .we_active(32'sd0),
  .num_byte_enables(32'sd1),
  .clock_edge(32'sd1),
  .no_of_RAM_readwrite_port(32'sd1)) mem_inst_banks_bank_array_impl_data6_rsc_comp
      (
      .data_in(mem_inst_banks_bank_array_impl_data6_rsc_data_in),
      .addr(mem_inst_banks_bank_array_impl_data6_rsc_addr),
      .re(mem_inst_banks_bank_array_impl_data6_rsc_re),
      .we(mem_inst_banks_bank_array_impl_data6_rsc_we),
      .data_out(mem_inst_banks_bank_array_impl_data6_rsc_data_out),
      .clk(clk),
      .a_rst(rst),
      .s_rst(1'b1),
      .en(mem_inst_banks_bank_array_impl_data6_rsc_en)
    );
  ram_sync_single_be #(.ram_id(32'sd304),
  .words(32'sd32),
  .width(32'sd8),
  .addr_width(32'sd5),
  .a_reset_active(32'sd0),
  .s_reset_active(32'sd0),
  .enable_active(32'sd0),
  .re_active(32'sd0),
  .we_active(32'sd0),
  .num_byte_enables(32'sd1),
  .clock_edge(32'sd1),
  .no_of_RAM_readwrite_port(32'sd1)) mem_inst_banks_bank_array_impl_data7_rsc_comp
      (
      .data_in(mem_inst_banks_bank_array_impl_data7_rsc_data_in),
      .addr(mem_inst_banks_bank_array_impl_data7_rsc_addr),
      .re(mem_inst_banks_bank_array_impl_data7_rsc_re),
      .we(mem_inst_banks_bank_array_impl_data7_rsc_we),
      .data_out(mem_inst_banks_bank_array_impl_data7_rsc_data_out),
      .clk(clk),
      .a_rst(rst),
      .s_rst(1'b1),
      .en(mem_inst_banks_bank_array_impl_data7_rsc_en)
    );
  InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_297_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
      mem_inst_banks_bank_array_impl_data0_rsci (
      .en(mem_inst_banks_bank_array_impl_data0_rsc_en),
      .data_out(mem_inst_banks_bank_array_impl_data0_rsc_data_out),
      .we(mem_inst_banks_bank_array_impl_data0_rsc_we),
      .re(mem_inst_banks_bank_array_impl_data0_rsc_re),
      .addr(mem_inst_banks_bank_array_impl_data0_rsc_addr),
      .data_in(mem_inst_banks_bank_array_impl_data0_rsc_data_in),
      .data_in_d(mem_inst_banks_bank_array_impl_data0_rsci_data_in_d),
      .addr_d(mem_inst_banks_bank_array_impl_data0_rsci_addr_d),
      .re_d(mem_inst_banks_bank_array_impl_data0_rsci_re_d),
      .we_d(mem_inst_banks_bank_array_impl_data0_rsci_we_d),
      .data_out_d(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d),
      .en_d(mem_inst_banks_bank_array_impl_data0_rsci_en_d)
    );
  InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_298_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
      mem_inst_banks_bank_array_impl_data1_rsci (
      .en(mem_inst_banks_bank_array_impl_data1_rsc_en),
      .data_out(mem_inst_banks_bank_array_impl_data1_rsc_data_out),
      .we(mem_inst_banks_bank_array_impl_data1_rsc_we),
      .re(mem_inst_banks_bank_array_impl_data1_rsc_re),
      .addr(mem_inst_banks_bank_array_impl_data1_rsc_addr),
      .data_in(mem_inst_banks_bank_array_impl_data1_rsc_data_in),
      .data_in_d(mem_inst_banks_bank_array_impl_data1_rsci_data_in_d),
      .addr_d(mem_inst_banks_bank_array_impl_data1_rsci_addr_d),
      .re_d(mem_inst_banks_bank_array_impl_data1_rsci_re_d),
      .we_d(mem_inst_banks_bank_array_impl_data1_rsci_we_d),
      .data_out_d(mem_inst_banks_bank_array_impl_data1_rsci_data_out_d),
      .en_d(mem_inst_banks_bank_array_impl_data1_rsci_en_d)
    );
  InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_299_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
      mem_inst_banks_bank_array_impl_data2_rsci (
      .en(mem_inst_banks_bank_array_impl_data2_rsc_en),
      .data_out(mem_inst_banks_bank_array_impl_data2_rsc_data_out),
      .we(mem_inst_banks_bank_array_impl_data2_rsc_we),
      .re(mem_inst_banks_bank_array_impl_data2_rsc_re),
      .addr(mem_inst_banks_bank_array_impl_data2_rsc_addr),
      .data_in(mem_inst_banks_bank_array_impl_data2_rsc_data_in),
      .data_in_d(mem_inst_banks_bank_array_impl_data2_rsci_data_in_d),
      .addr_d(mem_inst_banks_bank_array_impl_data2_rsci_addr_d),
      .re_d(mem_inst_banks_bank_array_impl_data2_rsci_re_d),
      .we_d(mem_inst_banks_bank_array_impl_data2_rsci_we_d),
      .data_out_d(mem_inst_banks_bank_array_impl_data2_rsci_data_out_d),
      .en_d(mem_inst_banks_bank_array_impl_data2_rsci_en_d)
    );
  InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_300_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
      mem_inst_banks_bank_array_impl_data3_rsci (
      .en(mem_inst_banks_bank_array_impl_data3_rsc_en),
      .data_out(mem_inst_banks_bank_array_impl_data3_rsc_data_out),
      .we(mem_inst_banks_bank_array_impl_data3_rsc_we),
      .re(mem_inst_banks_bank_array_impl_data3_rsc_re),
      .addr(mem_inst_banks_bank_array_impl_data3_rsc_addr),
      .data_in(mem_inst_banks_bank_array_impl_data3_rsc_data_in),
      .data_in_d(mem_inst_banks_bank_array_impl_data3_rsci_data_in_d),
      .addr_d(mem_inst_banks_bank_array_impl_data3_rsci_addr_d),
      .re_d(mem_inst_banks_bank_array_impl_data3_rsci_re_d),
      .we_d(mem_inst_banks_bank_array_impl_data3_rsci_we_d),
      .data_out_d(mem_inst_banks_bank_array_impl_data3_rsci_data_out_d),
      .en_d(mem_inst_banks_bank_array_impl_data3_rsci_en_d)
    );
  InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_301_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
      mem_inst_banks_bank_array_impl_data4_rsci (
      .en(mem_inst_banks_bank_array_impl_data4_rsc_en),
      .data_out(mem_inst_banks_bank_array_impl_data4_rsc_data_out),
      .we(mem_inst_banks_bank_array_impl_data4_rsc_we),
      .re(mem_inst_banks_bank_array_impl_data4_rsc_re),
      .addr(mem_inst_banks_bank_array_impl_data4_rsc_addr),
      .data_in(mem_inst_banks_bank_array_impl_data4_rsc_data_in),
      .data_in_d(mem_inst_banks_bank_array_impl_data4_rsci_data_in_d),
      .addr_d(mem_inst_banks_bank_array_impl_data4_rsci_addr_d),
      .re_d(mem_inst_banks_bank_array_impl_data4_rsci_re_d),
      .we_d(mem_inst_banks_bank_array_impl_data4_rsci_we_d),
      .data_out_d(mem_inst_banks_bank_array_impl_data4_rsci_data_out_d),
      .en_d(mem_inst_banks_bank_array_impl_data4_rsci_en_d)
    );
  InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_302_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
      mem_inst_banks_bank_array_impl_data5_rsci (
      .en(mem_inst_banks_bank_array_impl_data5_rsc_en),
      .data_out(mem_inst_banks_bank_array_impl_data5_rsc_data_out),
      .we(mem_inst_banks_bank_array_impl_data5_rsc_we),
      .re(mem_inst_banks_bank_array_impl_data5_rsc_re),
      .addr(mem_inst_banks_bank_array_impl_data5_rsc_addr),
      .data_in(mem_inst_banks_bank_array_impl_data5_rsc_data_in),
      .data_in_d(mem_inst_banks_bank_array_impl_data5_rsci_data_in_d),
      .addr_d(mem_inst_banks_bank_array_impl_data5_rsci_addr_d),
      .re_d(mem_inst_banks_bank_array_impl_data5_rsci_re_d),
      .we_d(mem_inst_banks_bank_array_impl_data5_rsci_we_d),
      .data_out_d(mem_inst_banks_bank_array_impl_data5_rsci_data_out_d),
      .en_d(mem_inst_banks_bank_array_impl_data5_rsci_en_d)
    );
  InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_303_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
      mem_inst_banks_bank_array_impl_data6_rsci (
      .en(mem_inst_banks_bank_array_impl_data6_rsc_en),
      .data_out(mem_inst_banks_bank_array_impl_data6_rsc_data_out),
      .we(mem_inst_banks_bank_array_impl_data6_rsc_we),
      .re(mem_inst_banks_bank_array_impl_data6_rsc_re),
      .addr(mem_inst_banks_bank_array_impl_data6_rsc_addr),
      .data_in(mem_inst_banks_bank_array_impl_data6_rsc_data_in),
      .data_in_d(mem_inst_banks_bank_array_impl_data6_rsci_data_in_d),
      .addr_d(mem_inst_banks_bank_array_impl_data6_rsci_addr_d),
      .re_d(mem_inst_banks_bank_array_impl_data6_rsci_re_d),
      .we_d(mem_inst_banks_bank_array_impl_data6_rsci_we_d),
      .data_out_d(mem_inst_banks_bank_array_impl_data6_rsci_data_out_d),
      .en_d(mem_inst_banks_bank_array_impl_data6_rsci_en_d)
    );
  InputSetup_ram_sample_065nm_singleport_beh_dc_RAM_rwport_en_304_32_8_5_0_0_0_0_0_1_1_32_8_1_gen
      mem_inst_banks_bank_array_impl_data7_rsci (
      .en(mem_inst_banks_bank_array_impl_data7_rsc_en),
      .data_out(mem_inst_banks_bank_array_impl_data7_rsc_data_out),
      .we(mem_inst_banks_bank_array_impl_data7_rsc_we),
      .re(mem_inst_banks_bank_array_impl_data7_rsc_re),
      .addr(mem_inst_banks_bank_array_impl_data7_rsc_addr),
      .data_in(mem_inst_banks_bank_array_impl_data7_rsc_data_in),
      .data_in_d(mem_inst_banks_bank_array_impl_data7_rsci_data_in_d),
      .addr_d(mem_inst_banks_bank_array_impl_data7_rsci_addr_d),
      .re_d(mem_inst_banks_bank_array_impl_data7_rsci_re_d),
      .we_d(mem_inst_banks_bank_array_impl_data7_rsci_we_d),
      .data_out_d(mem_inst_banks_bank_array_impl_data7_rsci_data_out_d),
      .en_d(mem_inst_banks_bank_array_impl_data7_rsci_en_d)
    );
  InputSetup_MemoryRun InputSetup_MemoryRun_inst (
      .clk(clk),
      .rst(rst),
      .write_req_val(write_req_val),
      .write_req_rdy(write_req_rdy),
      .write_req_msg(write_req_msg),
      .req_inter_val(req_inter_val),
      .req_inter_rdy(req_inter_rdy),
      .req_inter_msg(req_inter_msg),
      .rsp_inter_val(rsp_inter_val),
      .rsp_inter_rdy(rsp_inter_rdy),
      .rsp_inter_msg(rsp_inter_msg),
      .mem_inst_banks_bank_array_impl_data0_rsci_data_in_d(mem_inst_banks_bank_array_impl_data0_rsci_data_in_d),
      .mem_inst_banks_bank_array_impl_data0_rsci_addr_d(mem_inst_banks_bank_array_impl_data0_rsci_addr_d),
      .mem_inst_banks_bank_array_impl_data0_rsci_re_d(mem_inst_banks_bank_array_impl_data0_rsci_re_d),
      .mem_inst_banks_bank_array_impl_data0_rsci_we_d(mem_inst_banks_bank_array_impl_data0_rsci_we_d),
      .mem_inst_banks_bank_array_impl_data0_rsci_data_out_d(mem_inst_banks_bank_array_impl_data0_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data0_rsci_en_d(mem_inst_banks_bank_array_impl_data0_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data1_rsci_data_in_d(mem_inst_banks_bank_array_impl_data1_rsci_data_in_d),
      .mem_inst_banks_bank_array_impl_data1_rsci_addr_d(mem_inst_banks_bank_array_impl_data1_rsci_addr_d),
      .mem_inst_banks_bank_array_impl_data1_rsci_re_d(mem_inst_banks_bank_array_impl_data1_rsci_re_d),
      .mem_inst_banks_bank_array_impl_data1_rsci_we_d(mem_inst_banks_bank_array_impl_data1_rsci_we_d),
      .mem_inst_banks_bank_array_impl_data1_rsci_data_out_d(mem_inst_banks_bank_array_impl_data1_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data1_rsci_en_d(mem_inst_banks_bank_array_impl_data1_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data2_rsci_data_in_d(mem_inst_banks_bank_array_impl_data2_rsci_data_in_d),
      .mem_inst_banks_bank_array_impl_data2_rsci_addr_d(mem_inst_banks_bank_array_impl_data2_rsci_addr_d),
      .mem_inst_banks_bank_array_impl_data2_rsci_re_d(mem_inst_banks_bank_array_impl_data2_rsci_re_d),
      .mem_inst_banks_bank_array_impl_data2_rsci_we_d(mem_inst_banks_bank_array_impl_data2_rsci_we_d),
      .mem_inst_banks_bank_array_impl_data2_rsci_data_out_d(mem_inst_banks_bank_array_impl_data2_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data2_rsci_en_d(mem_inst_banks_bank_array_impl_data2_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data3_rsci_data_in_d(mem_inst_banks_bank_array_impl_data3_rsci_data_in_d),
      .mem_inst_banks_bank_array_impl_data3_rsci_addr_d(mem_inst_banks_bank_array_impl_data3_rsci_addr_d),
      .mem_inst_banks_bank_array_impl_data3_rsci_re_d(mem_inst_banks_bank_array_impl_data3_rsci_re_d),
      .mem_inst_banks_bank_array_impl_data3_rsci_we_d(mem_inst_banks_bank_array_impl_data3_rsci_we_d),
      .mem_inst_banks_bank_array_impl_data3_rsci_data_out_d(mem_inst_banks_bank_array_impl_data3_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data3_rsci_en_d(mem_inst_banks_bank_array_impl_data3_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data4_rsci_data_in_d(mem_inst_banks_bank_array_impl_data4_rsci_data_in_d),
      .mem_inst_banks_bank_array_impl_data4_rsci_addr_d(mem_inst_banks_bank_array_impl_data4_rsci_addr_d),
      .mem_inst_banks_bank_array_impl_data4_rsci_re_d(mem_inst_banks_bank_array_impl_data4_rsci_re_d),
      .mem_inst_banks_bank_array_impl_data4_rsci_we_d(mem_inst_banks_bank_array_impl_data4_rsci_we_d),
      .mem_inst_banks_bank_array_impl_data4_rsci_data_out_d(mem_inst_banks_bank_array_impl_data4_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data4_rsci_en_d(mem_inst_banks_bank_array_impl_data4_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data5_rsci_data_in_d(mem_inst_banks_bank_array_impl_data5_rsci_data_in_d),
      .mem_inst_banks_bank_array_impl_data5_rsci_addr_d(mem_inst_banks_bank_array_impl_data5_rsci_addr_d),
      .mem_inst_banks_bank_array_impl_data5_rsci_re_d(mem_inst_banks_bank_array_impl_data5_rsci_re_d),
      .mem_inst_banks_bank_array_impl_data5_rsci_we_d(mem_inst_banks_bank_array_impl_data5_rsci_we_d),
      .mem_inst_banks_bank_array_impl_data5_rsci_data_out_d(mem_inst_banks_bank_array_impl_data5_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data5_rsci_en_d(mem_inst_banks_bank_array_impl_data5_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data6_rsci_data_in_d(mem_inst_banks_bank_array_impl_data6_rsci_data_in_d),
      .mem_inst_banks_bank_array_impl_data6_rsci_addr_d(mem_inst_banks_bank_array_impl_data6_rsci_addr_d),
      .mem_inst_banks_bank_array_impl_data6_rsci_re_d(mem_inst_banks_bank_array_impl_data6_rsci_re_d),
      .mem_inst_banks_bank_array_impl_data6_rsci_we_d(mem_inst_banks_bank_array_impl_data6_rsci_we_d),
      .mem_inst_banks_bank_array_impl_data6_rsci_data_out_d(mem_inst_banks_bank_array_impl_data6_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data6_rsci_en_d(mem_inst_banks_bank_array_impl_data6_rsci_en_d),
      .mem_inst_banks_bank_array_impl_data7_rsci_data_in_d(mem_inst_banks_bank_array_impl_data7_rsci_data_in_d),
      .mem_inst_banks_bank_array_impl_data7_rsci_addr_d(mem_inst_banks_bank_array_impl_data7_rsci_addr_d),
      .mem_inst_banks_bank_array_impl_data7_rsci_re_d(mem_inst_banks_bank_array_impl_data7_rsci_re_d),
      .mem_inst_banks_bank_array_impl_data7_rsci_we_d(mem_inst_banks_bank_array_impl_data7_rsci_we_d),
      .mem_inst_banks_bank_array_impl_data7_rsci_data_out_d(mem_inst_banks_bank_array_impl_data7_rsci_data_out_d),
      .mem_inst_banks_bank_array_impl_data7_rsci_en_d(mem_inst_banks_bank_array_impl_data7_rsci_en_d)
    );
  InputSetup_ReadReqRun InputSetup_ReadReqRun_inst (
      .clk(clk),
      .rst(rst),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .req_inter_val(req_inter_val),
      .req_inter_rdy(req_inter_rdy),
      .req_inter_msg(req_inter_msg)
    );
  InputSetup_ReadRspRun InputSetup_ReadRspRun_inst (
      .clk(clk),
      .rst(rst),
      .act_in_vec_0_val(act_in_vec_0_val),
      .act_in_vec_1_val(act_in_vec_1_val),
      .act_in_vec_2_val(act_in_vec_2_val),
      .act_in_vec_3_val(act_in_vec_3_val),
      .act_in_vec_4_val(act_in_vec_4_val),
      .act_in_vec_5_val(act_in_vec_5_val),
      .act_in_vec_6_val(act_in_vec_6_val),
      .act_in_vec_7_val(act_in_vec_7_val),
      .act_in_vec_0_rdy(act_in_vec_0_rdy),
      .act_in_vec_1_rdy(act_in_vec_1_rdy),
      .act_in_vec_2_rdy(act_in_vec_2_rdy),
      .act_in_vec_3_rdy(act_in_vec_3_rdy),
      .act_in_vec_4_rdy(act_in_vec_4_rdy),
      .act_in_vec_5_rdy(act_in_vec_5_rdy),
      .act_in_vec_6_rdy(act_in_vec_6_rdy),
      .act_in_vec_7_rdy(act_in_vec_7_rdy),
      .act_in_vec_0_msg(act_in_vec_0_msg),
      .act_in_vec_1_msg(act_in_vec_1_msg),
      .act_in_vec_2_msg(act_in_vec_2_msg),
      .act_in_vec_3_msg(act_in_vec_3_msg),
      .act_in_vec_4_msg(act_in_vec_4_msg),
      .act_in_vec_5_msg(act_in_vec_5_msg),
      .act_in_vec_6_msg(act_in_vec_6_msg),
      .act_in_vec_7_msg(act_in_vec_7_msg),
      .rsp_inter_val(rsp_inter_val),
      .rsp_inter_rdy(rsp_inter_rdy),
      .rsp_inter_msg(rsp_inter_msg)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysArray
// ------------------------------------------------------------------


module SysArray (
  clk, rst, weight_in_vec_0_val, weight_in_vec_1_val, weight_in_vec_2_val, weight_in_vec_3_val,
      weight_in_vec_4_val, weight_in_vec_5_val, weight_in_vec_6_val, weight_in_vec_7_val,
      weight_in_vec_0_rdy, weight_in_vec_1_rdy, weight_in_vec_2_rdy, weight_in_vec_3_rdy,
      weight_in_vec_4_rdy, weight_in_vec_5_rdy, weight_in_vec_6_rdy, weight_in_vec_7_rdy,
      weight_in_vec_0_msg, weight_in_vec_1_msg, weight_in_vec_2_msg, weight_in_vec_3_msg,
      weight_in_vec_4_msg, weight_in_vec_5_msg, weight_in_vec_6_msg, weight_in_vec_7_msg,
      act_in_vec_0_val, act_in_vec_1_val, act_in_vec_2_val, act_in_vec_3_val, act_in_vec_4_val,
      act_in_vec_5_val, act_in_vec_6_val, act_in_vec_7_val, act_in_vec_0_rdy, act_in_vec_1_rdy,
      act_in_vec_2_rdy, act_in_vec_3_rdy, act_in_vec_4_rdy, act_in_vec_5_rdy, act_in_vec_6_rdy,
      act_in_vec_7_rdy, act_in_vec_0_msg, act_in_vec_1_msg, act_in_vec_2_msg, act_in_vec_3_msg,
      act_in_vec_4_msg, act_in_vec_5_msg, act_in_vec_6_msg, act_in_vec_7_msg, accum_out_vec_0_val,
      accum_out_vec_1_val, accum_out_vec_2_val, accum_out_vec_3_val, accum_out_vec_4_val,
      accum_out_vec_5_val, accum_out_vec_6_val, accum_out_vec_7_val, accum_out_vec_0_rdy,
      accum_out_vec_1_rdy, accum_out_vec_2_rdy, accum_out_vec_3_rdy, accum_out_vec_4_rdy,
      accum_out_vec_5_rdy, accum_out_vec_6_rdy, accum_out_vec_7_rdy, accum_out_vec_0_msg,
      accum_out_vec_1_msg, accum_out_vec_2_msg, accum_out_vec_3_msg, accum_out_vec_4_msg,
      accum_out_vec_5_msg, accum_out_vec_6_msg, accum_out_vec_7_msg
);
  input clk;
  input rst;
  input weight_in_vec_0_val;
  input weight_in_vec_1_val;
  input weight_in_vec_2_val;
  input weight_in_vec_3_val;
  input weight_in_vec_4_val;
  input weight_in_vec_5_val;
  input weight_in_vec_6_val;
  input weight_in_vec_7_val;
  output weight_in_vec_0_rdy;
  output weight_in_vec_1_rdy;
  output weight_in_vec_2_rdy;
  output weight_in_vec_3_rdy;
  output weight_in_vec_4_rdy;
  output weight_in_vec_5_rdy;
  output weight_in_vec_6_rdy;
  output weight_in_vec_7_rdy;
  input [7:0] weight_in_vec_0_msg;
  input [7:0] weight_in_vec_1_msg;
  input [7:0] weight_in_vec_2_msg;
  input [7:0] weight_in_vec_3_msg;
  input [7:0] weight_in_vec_4_msg;
  input [7:0] weight_in_vec_5_msg;
  input [7:0] weight_in_vec_6_msg;
  input [7:0] weight_in_vec_7_msg;
  input act_in_vec_0_val;
  input act_in_vec_1_val;
  input act_in_vec_2_val;
  input act_in_vec_3_val;
  input act_in_vec_4_val;
  input act_in_vec_5_val;
  input act_in_vec_6_val;
  input act_in_vec_7_val;
  output act_in_vec_0_rdy;
  output act_in_vec_1_rdy;
  output act_in_vec_2_rdy;
  output act_in_vec_3_rdy;
  output act_in_vec_4_rdy;
  output act_in_vec_5_rdy;
  output act_in_vec_6_rdy;
  output act_in_vec_7_rdy;
  input [7:0] act_in_vec_0_msg;
  input [7:0] act_in_vec_1_msg;
  input [7:0] act_in_vec_2_msg;
  input [7:0] act_in_vec_3_msg;
  input [7:0] act_in_vec_4_msg;
  input [7:0] act_in_vec_5_msg;
  input [7:0] act_in_vec_6_msg;
  input [7:0] act_in_vec_7_msg;
  output accum_out_vec_0_val;
  output accum_out_vec_1_val;
  output accum_out_vec_2_val;
  output accum_out_vec_3_val;
  output accum_out_vec_4_val;
  output accum_out_vec_5_val;
  output accum_out_vec_6_val;
  output accum_out_vec_7_val;
  input accum_out_vec_0_rdy;
  input accum_out_vec_1_rdy;
  input accum_out_vec_2_rdy;
  input accum_out_vec_3_rdy;
  input accum_out_vec_4_rdy;
  input accum_out_vec_5_rdy;
  input accum_out_vec_6_rdy;
  input accum_out_vec_7_rdy;
  output [31:0] accum_out_vec_0_msg;
  output [31:0] accum_out_vec_1_msg;
  output [31:0] accum_out_vec_2_msg;
  output [31:0] accum_out_vec_3_msg;
  output [31:0] accum_out_vec_4_msg;
  output [31:0] accum_out_vec_5_msg;
  output [31:0] accum_out_vec_6_msg;
  output [31:0] accum_out_vec_7_msg;


  // Interconnect Declarations
  wire weight_inter_0_0_val;
  wire weight_inter_0_1_val;
  wire weight_inter_0_2_val;
  wire weight_inter_0_3_val;
  wire weight_inter_0_4_val;
  wire weight_inter_0_5_val;
  wire weight_inter_0_6_val;
  wire weight_inter_0_7_val;
  wire weight_inter_1_0_val;
  wire weight_inter_1_1_val;
  wire weight_inter_1_2_val;
  wire weight_inter_1_3_val;
  wire weight_inter_1_4_val;
  wire weight_inter_1_5_val;
  wire weight_inter_1_6_val;
  wire weight_inter_1_7_val;
  wire weight_inter_2_0_val;
  wire weight_inter_2_1_val;
  wire weight_inter_2_2_val;
  wire weight_inter_2_3_val;
  wire weight_inter_2_4_val;
  wire weight_inter_2_5_val;
  wire weight_inter_2_6_val;
  wire weight_inter_2_7_val;
  wire weight_inter_3_0_val;
  wire weight_inter_3_1_val;
  wire weight_inter_3_2_val;
  wire weight_inter_3_3_val;
  wire weight_inter_3_4_val;
  wire weight_inter_3_5_val;
  wire weight_inter_3_6_val;
  wire weight_inter_3_7_val;
  wire weight_inter_4_0_val;
  wire weight_inter_4_1_val;
  wire weight_inter_4_2_val;
  wire weight_inter_4_3_val;
  wire weight_inter_4_4_val;
  wire weight_inter_4_5_val;
  wire weight_inter_4_6_val;
  wire weight_inter_4_7_val;
  wire weight_inter_5_0_val;
  wire weight_inter_5_1_val;
  wire weight_inter_5_2_val;
  wire weight_inter_5_3_val;
  wire weight_inter_5_4_val;
  wire weight_inter_5_5_val;
  wire weight_inter_5_6_val;
  wire weight_inter_5_7_val;
  wire weight_inter_6_0_val;
  wire weight_inter_6_1_val;
  wire weight_inter_6_2_val;
  wire weight_inter_6_3_val;
  wire weight_inter_6_4_val;
  wire weight_inter_6_5_val;
  wire weight_inter_6_6_val;
  wire weight_inter_6_7_val;
  wire weight_inter_7_0_val;
  wire weight_inter_7_1_val;
  wire weight_inter_7_2_val;
  wire weight_inter_7_3_val;
  wire weight_inter_7_4_val;
  wire weight_inter_7_5_val;
  wire weight_inter_7_6_val;
  wire weight_inter_7_7_val;
  wire weight_inter_0_0_rdy;
  wire weight_inter_0_1_rdy;
  wire weight_inter_0_2_rdy;
  wire weight_inter_0_3_rdy;
  wire weight_inter_0_4_rdy;
  wire weight_inter_0_5_rdy;
  wire weight_inter_0_6_rdy;
  wire weight_inter_0_7_rdy;
  wire weight_inter_1_0_rdy;
  wire weight_inter_1_1_rdy;
  wire weight_inter_1_2_rdy;
  wire weight_inter_1_3_rdy;
  wire weight_inter_1_4_rdy;
  wire weight_inter_1_5_rdy;
  wire weight_inter_1_6_rdy;
  wire weight_inter_1_7_rdy;
  wire weight_inter_2_0_rdy;
  wire weight_inter_2_1_rdy;
  wire weight_inter_2_2_rdy;
  wire weight_inter_2_3_rdy;
  wire weight_inter_2_4_rdy;
  wire weight_inter_2_5_rdy;
  wire weight_inter_2_6_rdy;
  wire weight_inter_2_7_rdy;
  wire weight_inter_3_0_rdy;
  wire weight_inter_3_1_rdy;
  wire weight_inter_3_2_rdy;
  wire weight_inter_3_3_rdy;
  wire weight_inter_3_4_rdy;
  wire weight_inter_3_5_rdy;
  wire weight_inter_3_6_rdy;
  wire weight_inter_3_7_rdy;
  wire weight_inter_4_0_rdy;
  wire weight_inter_4_1_rdy;
  wire weight_inter_4_2_rdy;
  wire weight_inter_4_3_rdy;
  wire weight_inter_4_4_rdy;
  wire weight_inter_4_5_rdy;
  wire weight_inter_4_6_rdy;
  wire weight_inter_4_7_rdy;
  wire weight_inter_5_0_rdy;
  wire weight_inter_5_1_rdy;
  wire weight_inter_5_2_rdy;
  wire weight_inter_5_3_rdy;
  wire weight_inter_5_4_rdy;
  wire weight_inter_5_5_rdy;
  wire weight_inter_5_6_rdy;
  wire weight_inter_5_7_rdy;
  wire weight_inter_6_0_rdy;
  wire weight_inter_6_1_rdy;
  wire weight_inter_6_2_rdy;
  wire weight_inter_6_3_rdy;
  wire weight_inter_6_4_rdy;
  wire weight_inter_6_5_rdy;
  wire weight_inter_6_6_rdy;
  wire weight_inter_6_7_rdy;
  wire weight_inter_7_0_rdy;
  wire weight_inter_7_1_rdy;
  wire weight_inter_7_2_rdy;
  wire weight_inter_7_3_rdy;
  wire weight_inter_7_4_rdy;
  wire weight_inter_7_5_rdy;
  wire weight_inter_7_6_rdy;
  wire weight_inter_7_7_rdy;
  wire [7:0] weight_inter_0_0_msg;
  wire [7:0] weight_inter_0_1_msg;
  wire [7:0] weight_inter_0_2_msg;
  wire [7:0] weight_inter_0_3_msg;
  wire [7:0] weight_inter_0_4_msg;
  wire [7:0] weight_inter_0_5_msg;
  wire [7:0] weight_inter_0_6_msg;
  wire [7:0] weight_inter_0_7_msg;
  wire [7:0] weight_inter_1_0_msg;
  wire [7:0] weight_inter_1_1_msg;
  wire [7:0] weight_inter_1_2_msg;
  wire [7:0] weight_inter_1_3_msg;
  wire [7:0] weight_inter_1_4_msg;
  wire [7:0] weight_inter_1_5_msg;
  wire [7:0] weight_inter_1_6_msg;
  wire [7:0] weight_inter_1_7_msg;
  wire [7:0] weight_inter_2_0_msg;
  wire [7:0] weight_inter_2_1_msg;
  wire [7:0] weight_inter_2_2_msg;
  wire [7:0] weight_inter_2_3_msg;
  wire [7:0] weight_inter_2_4_msg;
  wire [7:0] weight_inter_2_5_msg;
  wire [7:0] weight_inter_2_6_msg;
  wire [7:0] weight_inter_2_7_msg;
  wire [7:0] weight_inter_3_0_msg;
  wire [7:0] weight_inter_3_1_msg;
  wire [7:0] weight_inter_3_2_msg;
  wire [7:0] weight_inter_3_3_msg;
  wire [7:0] weight_inter_3_4_msg;
  wire [7:0] weight_inter_3_5_msg;
  wire [7:0] weight_inter_3_6_msg;
  wire [7:0] weight_inter_3_7_msg;
  wire [7:0] weight_inter_4_0_msg;
  wire [7:0] weight_inter_4_1_msg;
  wire [7:0] weight_inter_4_2_msg;
  wire [7:0] weight_inter_4_3_msg;
  wire [7:0] weight_inter_4_4_msg;
  wire [7:0] weight_inter_4_5_msg;
  wire [7:0] weight_inter_4_6_msg;
  wire [7:0] weight_inter_4_7_msg;
  wire [7:0] weight_inter_5_0_msg;
  wire [7:0] weight_inter_5_1_msg;
  wire [7:0] weight_inter_5_2_msg;
  wire [7:0] weight_inter_5_3_msg;
  wire [7:0] weight_inter_5_4_msg;
  wire [7:0] weight_inter_5_5_msg;
  wire [7:0] weight_inter_5_6_msg;
  wire [7:0] weight_inter_5_7_msg;
  wire [7:0] weight_inter_6_0_msg;
  wire [7:0] weight_inter_6_1_msg;
  wire [7:0] weight_inter_6_2_msg;
  wire [7:0] weight_inter_6_3_msg;
  wire [7:0] weight_inter_6_4_msg;
  wire [7:0] weight_inter_6_5_msg;
  wire [7:0] weight_inter_6_6_msg;
  wire [7:0] weight_inter_6_7_msg;
  wire [7:0] weight_inter_7_0_msg;
  wire [7:0] weight_inter_7_1_msg;
  wire [7:0] weight_inter_7_2_msg;
  wire [7:0] weight_inter_7_3_msg;
  wire [7:0] weight_inter_7_4_msg;
  wire [7:0] weight_inter_7_5_msg;
  wire [7:0] weight_inter_7_6_msg;
  wire [7:0] weight_inter_7_7_msg;
  wire act_inter_0_0_val;
  wire act_inter_0_1_val;
  wire act_inter_0_2_val;
  wire act_inter_0_3_val;
  wire act_inter_0_4_val;
  wire act_inter_0_5_val;
  wire act_inter_0_6_val;
  wire act_inter_0_7_val;
  wire act_inter_1_0_val;
  wire act_inter_1_1_val;
  wire act_inter_1_2_val;
  wire act_inter_1_3_val;
  wire act_inter_1_4_val;
  wire act_inter_1_5_val;
  wire act_inter_1_6_val;
  wire act_inter_1_7_val;
  wire act_inter_2_0_val;
  wire act_inter_2_1_val;
  wire act_inter_2_2_val;
  wire act_inter_2_3_val;
  wire act_inter_2_4_val;
  wire act_inter_2_5_val;
  wire act_inter_2_6_val;
  wire act_inter_2_7_val;
  wire act_inter_3_0_val;
  wire act_inter_3_1_val;
  wire act_inter_3_2_val;
  wire act_inter_3_3_val;
  wire act_inter_3_4_val;
  wire act_inter_3_5_val;
  wire act_inter_3_6_val;
  wire act_inter_3_7_val;
  wire act_inter_4_0_val;
  wire act_inter_4_1_val;
  wire act_inter_4_2_val;
  wire act_inter_4_3_val;
  wire act_inter_4_4_val;
  wire act_inter_4_5_val;
  wire act_inter_4_6_val;
  wire act_inter_4_7_val;
  wire act_inter_5_0_val;
  wire act_inter_5_1_val;
  wire act_inter_5_2_val;
  wire act_inter_5_3_val;
  wire act_inter_5_4_val;
  wire act_inter_5_5_val;
  wire act_inter_5_6_val;
  wire act_inter_5_7_val;
  wire act_inter_6_0_val;
  wire act_inter_6_1_val;
  wire act_inter_6_2_val;
  wire act_inter_6_3_val;
  wire act_inter_6_4_val;
  wire act_inter_6_5_val;
  wire act_inter_6_6_val;
  wire act_inter_6_7_val;
  wire act_inter_7_0_val;
  wire act_inter_7_1_val;
  wire act_inter_7_2_val;
  wire act_inter_7_3_val;
  wire act_inter_7_4_val;
  wire act_inter_7_5_val;
  wire act_inter_7_6_val;
  wire act_inter_7_7_val;
  wire act_inter_0_0_rdy;
  wire act_inter_0_1_rdy;
  wire act_inter_0_2_rdy;
  wire act_inter_0_3_rdy;
  wire act_inter_0_4_rdy;
  wire act_inter_0_5_rdy;
  wire act_inter_0_6_rdy;
  wire act_inter_0_7_rdy;
  wire act_inter_1_0_rdy;
  wire act_inter_1_1_rdy;
  wire act_inter_1_2_rdy;
  wire act_inter_1_3_rdy;
  wire act_inter_1_4_rdy;
  wire act_inter_1_5_rdy;
  wire act_inter_1_6_rdy;
  wire act_inter_1_7_rdy;
  wire act_inter_2_0_rdy;
  wire act_inter_2_1_rdy;
  wire act_inter_2_2_rdy;
  wire act_inter_2_3_rdy;
  wire act_inter_2_4_rdy;
  wire act_inter_2_5_rdy;
  wire act_inter_2_6_rdy;
  wire act_inter_2_7_rdy;
  wire act_inter_3_0_rdy;
  wire act_inter_3_1_rdy;
  wire act_inter_3_2_rdy;
  wire act_inter_3_3_rdy;
  wire act_inter_3_4_rdy;
  wire act_inter_3_5_rdy;
  wire act_inter_3_6_rdy;
  wire act_inter_3_7_rdy;
  wire act_inter_4_0_rdy;
  wire act_inter_4_1_rdy;
  wire act_inter_4_2_rdy;
  wire act_inter_4_3_rdy;
  wire act_inter_4_4_rdy;
  wire act_inter_4_5_rdy;
  wire act_inter_4_6_rdy;
  wire act_inter_4_7_rdy;
  wire act_inter_5_0_rdy;
  wire act_inter_5_1_rdy;
  wire act_inter_5_2_rdy;
  wire act_inter_5_3_rdy;
  wire act_inter_5_4_rdy;
  wire act_inter_5_5_rdy;
  wire act_inter_5_6_rdy;
  wire act_inter_5_7_rdy;
  wire act_inter_6_0_rdy;
  wire act_inter_6_1_rdy;
  wire act_inter_6_2_rdy;
  wire act_inter_6_3_rdy;
  wire act_inter_6_4_rdy;
  wire act_inter_6_5_rdy;
  wire act_inter_6_6_rdy;
  wire act_inter_6_7_rdy;
  wire act_inter_7_0_rdy;
  wire act_inter_7_1_rdy;
  wire act_inter_7_2_rdy;
  wire act_inter_7_3_rdy;
  wire act_inter_7_4_rdy;
  wire act_inter_7_5_rdy;
  wire act_inter_7_6_rdy;
  wire act_inter_7_7_rdy;
  wire [7:0] act_inter_0_0_msg;
  wire [7:0] act_inter_0_1_msg;
  wire [7:0] act_inter_0_2_msg;
  wire [7:0] act_inter_0_3_msg;
  wire [7:0] act_inter_0_4_msg;
  wire [7:0] act_inter_0_5_msg;
  wire [7:0] act_inter_0_6_msg;
  wire [7:0] act_inter_0_7_msg;
  wire [7:0] act_inter_1_0_msg;
  wire [7:0] act_inter_1_1_msg;
  wire [7:0] act_inter_1_2_msg;
  wire [7:0] act_inter_1_3_msg;
  wire [7:0] act_inter_1_4_msg;
  wire [7:0] act_inter_1_5_msg;
  wire [7:0] act_inter_1_6_msg;
  wire [7:0] act_inter_1_7_msg;
  wire [7:0] act_inter_2_0_msg;
  wire [7:0] act_inter_2_1_msg;
  wire [7:0] act_inter_2_2_msg;
  wire [7:0] act_inter_2_3_msg;
  wire [7:0] act_inter_2_4_msg;
  wire [7:0] act_inter_2_5_msg;
  wire [7:0] act_inter_2_6_msg;
  wire [7:0] act_inter_2_7_msg;
  wire [7:0] act_inter_3_0_msg;
  wire [7:0] act_inter_3_1_msg;
  wire [7:0] act_inter_3_2_msg;
  wire [7:0] act_inter_3_3_msg;
  wire [7:0] act_inter_3_4_msg;
  wire [7:0] act_inter_3_5_msg;
  wire [7:0] act_inter_3_6_msg;
  wire [7:0] act_inter_3_7_msg;
  wire [7:0] act_inter_4_0_msg;
  wire [7:0] act_inter_4_1_msg;
  wire [7:0] act_inter_4_2_msg;
  wire [7:0] act_inter_4_3_msg;
  wire [7:0] act_inter_4_4_msg;
  wire [7:0] act_inter_4_5_msg;
  wire [7:0] act_inter_4_6_msg;
  wire [7:0] act_inter_4_7_msg;
  wire [7:0] act_inter_5_0_msg;
  wire [7:0] act_inter_5_1_msg;
  wire [7:0] act_inter_5_2_msg;
  wire [7:0] act_inter_5_3_msg;
  wire [7:0] act_inter_5_4_msg;
  wire [7:0] act_inter_5_5_msg;
  wire [7:0] act_inter_5_6_msg;
  wire [7:0] act_inter_5_7_msg;
  wire [7:0] act_inter_6_0_msg;
  wire [7:0] act_inter_6_1_msg;
  wire [7:0] act_inter_6_2_msg;
  wire [7:0] act_inter_6_3_msg;
  wire [7:0] act_inter_6_4_msg;
  wire [7:0] act_inter_6_5_msg;
  wire [7:0] act_inter_6_6_msg;
  wire [7:0] act_inter_6_7_msg;
  wire [7:0] act_inter_7_0_msg;
  wire [7:0] act_inter_7_1_msg;
  wire [7:0] act_inter_7_2_msg;
  wire [7:0] act_inter_7_3_msg;
  wire [7:0] act_inter_7_4_msg;
  wire [7:0] act_inter_7_5_msg;
  wire [7:0] act_inter_7_6_msg;
  wire [7:0] act_inter_7_7_msg;
  wire accum_inter_0_0_val;
  wire accum_inter_0_1_val;
  wire accum_inter_0_2_val;
  wire accum_inter_0_3_val;
  wire accum_inter_0_4_val;
  wire accum_inter_0_5_val;
  wire accum_inter_0_6_val;
  wire accum_inter_0_7_val;
  wire accum_inter_1_0_val;
  wire accum_inter_1_1_val;
  wire accum_inter_1_2_val;
  wire accum_inter_1_3_val;
  wire accum_inter_1_4_val;
  wire accum_inter_1_5_val;
  wire accum_inter_1_6_val;
  wire accum_inter_1_7_val;
  wire accum_inter_2_0_val;
  wire accum_inter_2_1_val;
  wire accum_inter_2_2_val;
  wire accum_inter_2_3_val;
  wire accum_inter_2_4_val;
  wire accum_inter_2_5_val;
  wire accum_inter_2_6_val;
  wire accum_inter_2_7_val;
  wire accum_inter_3_0_val;
  wire accum_inter_3_1_val;
  wire accum_inter_3_2_val;
  wire accum_inter_3_3_val;
  wire accum_inter_3_4_val;
  wire accum_inter_3_5_val;
  wire accum_inter_3_6_val;
  wire accum_inter_3_7_val;
  wire accum_inter_4_0_val;
  wire accum_inter_4_1_val;
  wire accum_inter_4_2_val;
  wire accum_inter_4_3_val;
  wire accum_inter_4_4_val;
  wire accum_inter_4_5_val;
  wire accum_inter_4_6_val;
  wire accum_inter_4_7_val;
  wire accum_inter_5_0_val;
  wire accum_inter_5_1_val;
  wire accum_inter_5_2_val;
  wire accum_inter_5_3_val;
  wire accum_inter_5_4_val;
  wire accum_inter_5_5_val;
  wire accum_inter_5_6_val;
  wire accum_inter_5_7_val;
  wire accum_inter_6_0_val;
  wire accum_inter_6_1_val;
  wire accum_inter_6_2_val;
  wire accum_inter_6_3_val;
  wire accum_inter_6_4_val;
  wire accum_inter_6_5_val;
  wire accum_inter_6_6_val;
  wire accum_inter_6_7_val;
  wire accum_inter_7_0_val;
  wire accum_inter_7_1_val;
  wire accum_inter_7_2_val;
  wire accum_inter_7_3_val;
  wire accum_inter_7_4_val;
  wire accum_inter_7_5_val;
  wire accum_inter_7_6_val;
  wire accum_inter_7_7_val;
  wire accum_inter_0_0_rdy;
  wire accum_inter_0_1_rdy;
  wire accum_inter_0_2_rdy;
  wire accum_inter_0_3_rdy;
  wire accum_inter_0_4_rdy;
  wire accum_inter_0_5_rdy;
  wire accum_inter_0_6_rdy;
  wire accum_inter_0_7_rdy;
  wire accum_inter_1_0_rdy;
  wire accum_inter_1_1_rdy;
  wire accum_inter_1_2_rdy;
  wire accum_inter_1_3_rdy;
  wire accum_inter_1_4_rdy;
  wire accum_inter_1_5_rdy;
  wire accum_inter_1_6_rdy;
  wire accum_inter_1_7_rdy;
  wire accum_inter_2_0_rdy;
  wire accum_inter_2_1_rdy;
  wire accum_inter_2_2_rdy;
  wire accum_inter_2_3_rdy;
  wire accum_inter_2_4_rdy;
  wire accum_inter_2_5_rdy;
  wire accum_inter_2_6_rdy;
  wire accum_inter_2_7_rdy;
  wire accum_inter_3_0_rdy;
  wire accum_inter_3_1_rdy;
  wire accum_inter_3_2_rdy;
  wire accum_inter_3_3_rdy;
  wire accum_inter_3_4_rdy;
  wire accum_inter_3_5_rdy;
  wire accum_inter_3_6_rdy;
  wire accum_inter_3_7_rdy;
  wire accum_inter_4_0_rdy;
  wire accum_inter_4_1_rdy;
  wire accum_inter_4_2_rdy;
  wire accum_inter_4_3_rdy;
  wire accum_inter_4_4_rdy;
  wire accum_inter_4_5_rdy;
  wire accum_inter_4_6_rdy;
  wire accum_inter_4_7_rdy;
  wire accum_inter_5_0_rdy;
  wire accum_inter_5_1_rdy;
  wire accum_inter_5_2_rdy;
  wire accum_inter_5_3_rdy;
  wire accum_inter_5_4_rdy;
  wire accum_inter_5_5_rdy;
  wire accum_inter_5_6_rdy;
  wire accum_inter_5_7_rdy;
  wire accum_inter_6_0_rdy;
  wire accum_inter_6_1_rdy;
  wire accum_inter_6_2_rdy;
  wire accum_inter_6_3_rdy;
  wire accum_inter_6_4_rdy;
  wire accum_inter_6_5_rdy;
  wire accum_inter_6_6_rdy;
  wire accum_inter_6_7_rdy;
  wire accum_inter_7_0_rdy;
  wire accum_inter_7_1_rdy;
  wire accum_inter_7_2_rdy;
  wire accum_inter_7_3_rdy;
  wire accum_inter_7_4_rdy;
  wire accum_inter_7_5_rdy;
  wire accum_inter_7_6_rdy;
  wire accum_inter_7_7_rdy;
  wire [31:0] accum_inter_0_0_msg;
  wire [31:0] accum_inter_0_1_msg;
  wire [31:0] accum_inter_0_2_msg;
  wire [31:0] accum_inter_0_3_msg;
  wire [31:0] accum_inter_0_4_msg;
  wire [31:0] accum_inter_0_5_msg;
  wire [31:0] accum_inter_0_6_msg;
  wire [31:0] accum_inter_0_7_msg;
  wire [31:0] accum_inter_1_0_msg;
  wire [31:0] accum_inter_1_1_msg;
  wire [31:0] accum_inter_1_2_msg;
  wire [31:0] accum_inter_1_3_msg;
  wire [31:0] accum_inter_1_4_msg;
  wire [31:0] accum_inter_1_5_msg;
  wire [31:0] accum_inter_1_6_msg;
  wire [31:0] accum_inter_1_7_msg;
  wire [31:0] accum_inter_2_0_msg;
  wire [31:0] accum_inter_2_1_msg;
  wire [31:0] accum_inter_2_2_msg;
  wire [31:0] accum_inter_2_3_msg;
  wire [31:0] accum_inter_2_4_msg;
  wire [31:0] accum_inter_2_5_msg;
  wire [31:0] accum_inter_2_6_msg;
  wire [31:0] accum_inter_2_7_msg;
  wire [31:0] accum_inter_3_0_msg;
  wire [31:0] accum_inter_3_1_msg;
  wire [31:0] accum_inter_3_2_msg;
  wire [31:0] accum_inter_3_3_msg;
  wire [31:0] accum_inter_3_4_msg;
  wire [31:0] accum_inter_3_5_msg;
  wire [31:0] accum_inter_3_6_msg;
  wire [31:0] accum_inter_3_7_msg;
  wire [31:0] accum_inter_4_0_msg;
  wire [31:0] accum_inter_4_1_msg;
  wire [31:0] accum_inter_4_2_msg;
  wire [31:0] accum_inter_4_3_msg;
  wire [31:0] accum_inter_4_4_msg;
  wire [31:0] accum_inter_4_5_msg;
  wire [31:0] accum_inter_4_6_msg;
  wire [31:0] accum_inter_4_7_msg;
  wire [31:0] accum_inter_5_0_msg;
  wire [31:0] accum_inter_5_1_msg;
  wire [31:0] accum_inter_5_2_msg;
  wire [31:0] accum_inter_5_3_msg;
  wire [31:0] accum_inter_5_4_msg;
  wire [31:0] accum_inter_5_5_msg;
  wire [31:0] accum_inter_5_6_msg;
  wire [31:0] accum_inter_5_7_msg;
  wire [31:0] accum_inter_6_0_msg;
  wire [31:0] accum_inter_6_1_msg;
  wire [31:0] accum_inter_6_2_msg;
  wire [31:0] accum_inter_6_3_msg;
  wire [31:0] accum_inter_6_4_msg;
  wire [31:0] accum_inter_6_5_msg;
  wire [31:0] accum_inter_6_6_msg;
  wire [31:0] accum_inter_6_7_msg;
  wire [31:0] accum_inter_7_0_msg;
  wire [31:0] accum_inter_7_1_msg;
  wire [31:0] accum_inter_7_2_msg;
  wire [31:0] accum_inter_7_3_msg;
  wire [31:0] accum_inter_7_4_msg;
  wire [31:0] accum_inter_7_5_msg;
  wire [31:0] accum_inter_7_6_msg;
  wire [31:0] accum_inter_7_7_msg;
  wire [7:0] weight_inter_PopNB_56_mioi_data_rsc_z;
  wire weight_inter_PopNB_56_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_57_mioi_data_rsc_z;
  wire weight_inter_PopNB_57_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_58_mioi_data_rsc_z;
  wire weight_inter_PopNB_58_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_59_mioi_data_rsc_z;
  wire weight_inter_PopNB_59_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_60_mioi_data_rsc_z;
  wire weight_inter_PopNB_60_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_61_mioi_data_rsc_z;
  wire weight_inter_PopNB_61_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_62_mioi_data_rsc_z;
  wire weight_inter_PopNB_62_mioi_return_rsc_z;
  wire [7:0] weight_inter_PopNB_63_mioi_data_rsc_z;
  wire weight_inter_PopNB_63_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_7_mioi_data_rsc_z;
  wire act_inter_PopNB_7_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_15_mioi_data_rsc_z;
  wire act_inter_PopNB_15_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_23_mioi_data_rsc_z;
  wire act_inter_PopNB_23_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_31_mioi_data_rsc_z;
  wire act_inter_PopNB_31_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_39_mioi_data_rsc_z;
  wire act_inter_PopNB_39_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_47_mioi_data_rsc_z;
  wire act_inter_PopNB_47_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_55_mioi_data_rsc_z;
  wire act_inter_PopNB_55_mioi_return_rsc_z;
  wire [7:0] act_inter_PopNB_63_mioi_data_rsc_z;
  wire act_inter_PopNB_63_mioi_return_rsc_z;
  wire accum_inter_PushNB_mioi_return_rsc_z;
  wire accum_inter_PushNB_1_mioi_return_rsc_z;
  wire accum_inter_PushNB_2_mioi_return_rsc_z;
  wire accum_inter_PushNB_3_mioi_return_rsc_z;
  wire accum_inter_PushNB_4_mioi_return_rsc_z;
  wire accum_inter_PushNB_5_mioi_return_rsc_z;
  wire accum_inter_PushNB_6_mioi_return_rsc_z;
  wire accum_inter_PushNB_7_mioi_return_rsc_z;
  wire weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff;
  wire act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff;
  wire accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff;


  // Interconnect Declarations for Component Instantiations 
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_56_mioi
      (
      .this_val(weight_inter_7_0_val),
      .this_rdy(weight_inter_7_0_rdy),
      .this_msg(weight_inter_7_0_msg),
      .data_rsc_z(weight_inter_PopNB_56_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_56_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_57_mioi
      (
      .this_val(weight_inter_7_1_val),
      .this_rdy(weight_inter_7_1_rdy),
      .this_msg(weight_inter_7_1_msg),
      .data_rsc_z(weight_inter_PopNB_57_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_57_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_58_mioi
      (
      .this_val(weight_inter_7_2_val),
      .this_rdy(weight_inter_7_2_rdy),
      .this_msg(weight_inter_7_2_msg),
      .data_rsc_z(weight_inter_PopNB_58_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_58_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_59_mioi
      (
      .this_val(weight_inter_7_3_val),
      .this_rdy(weight_inter_7_3_rdy),
      .this_msg(weight_inter_7_3_msg),
      .data_rsc_z(weight_inter_PopNB_59_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_59_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_60_mioi
      (
      .this_val(weight_inter_7_4_val),
      .this_rdy(weight_inter_7_4_rdy),
      .this_msg(weight_inter_7_4_msg),
      .data_rsc_z(weight_inter_PopNB_60_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_60_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_61_mioi
      (
      .this_val(weight_inter_7_5_val),
      .this_rdy(weight_inter_7_5_rdy),
      .this_msg(weight_inter_7_5_msg),
      .data_rsc_z(weight_inter_PopNB_61_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_61_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_62_mioi
      (
      .this_val(weight_inter_7_6_val),
      .this_rdy(weight_inter_7_6_rdy),
      .this_msg(weight_inter_7_6_msg),
      .data_rsc_z(weight_inter_PopNB_62_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_62_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  weight_inter_PopNB_63_mioi
      (
      .this_val(weight_inter_7_7_val),
      .this_rdy(weight_inter_7_7_rdy),
      .this_msg(weight_inter_7_7_msg),
      .data_rsc_z(weight_inter_PopNB_63_mioi_data_rsc_z),
      .return_rsc_z(weight_inter_PopNB_63_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_7_mioi
      (
      .this_val(act_inter_0_7_val),
      .this_rdy(act_inter_0_7_rdy),
      .this_msg(act_inter_0_7_msg),
      .data_rsc_z(act_inter_PopNB_7_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_7_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_15_mioi
      (
      .this_val(act_inter_1_7_val),
      .this_rdy(act_inter_1_7_rdy),
      .this_msg(act_inter_1_7_msg),
      .data_rsc_z(act_inter_PopNB_15_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_15_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_23_mioi
      (
      .this_val(act_inter_2_7_val),
      .this_rdy(act_inter_2_7_rdy),
      .this_msg(act_inter_2_7_msg),
      .data_rsc_z(act_inter_PopNB_23_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_23_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_31_mioi
      (
      .this_val(act_inter_3_7_val),
      .this_rdy(act_inter_3_7_rdy),
      .this_msg(act_inter_3_7_msg),
      .data_rsc_z(act_inter_PopNB_31_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_31_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_39_mioi
      (
      .this_val(act_inter_4_7_val),
      .this_rdy(act_inter_4_7_rdy),
      .this_msg(act_inter_4_7_msg),
      .data_rsc_z(act_inter_PopNB_39_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_39_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_47_mioi
      (
      .this_val(act_inter_5_7_val),
      .this_rdy(act_inter_5_7_rdy),
      .this_msg(act_inter_5_7_msg),
      .data_rsc_z(act_inter_PopNB_47_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_47_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_55_mioi
      (
      .this_val(act_inter_6_7_val),
      .this_rdy(act_inter_6_7_rdy),
      .this_msg(act_inter_6_7_msg),
      .data_rsc_z(act_inter_PopNB_55_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_55_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_InputType_Connections_SYN_PORT_PopNB  act_inter_PopNB_63_mioi
      (
      .this_val(act_inter_7_7_val),
      .this_rdy(act_inter_7_7_rdy),
      .this_msg(act_inter_7_7_msg),
      .data_rsc_z(act_inter_PopNB_63_mioi_data_rsc_z),
      .return_rsc_z(act_inter_PopNB_63_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_mioi
      (
      .this_val(accum_inter_0_0_val),
      .this_rdy(accum_inter_0_0_rdy),
      .this_msg(accum_inter_0_0_msg),
      .return_rsc_z(accum_inter_PushNB_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_1_mioi
      (
      .this_val(accum_inter_0_1_val),
      .this_rdy(accum_inter_0_1_rdy),
      .this_msg(accum_inter_0_1_msg),
      .return_rsc_z(accum_inter_PushNB_1_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_2_mioi
      (
      .this_val(accum_inter_0_2_val),
      .this_rdy(accum_inter_0_2_rdy),
      .this_msg(accum_inter_0_2_msg),
      .return_rsc_z(accum_inter_PushNB_2_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_3_mioi
      (
      .this_val(accum_inter_0_3_val),
      .this_rdy(accum_inter_0_3_rdy),
      .this_msg(accum_inter_0_3_msg),
      .return_rsc_z(accum_inter_PushNB_3_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_4_mioi
      (
      .this_val(accum_inter_0_4_val),
      .this_rdy(accum_inter_0_4_rdy),
      .this_msg(accum_inter_0_4_msg),
      .return_rsc_z(accum_inter_PushNB_4_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_5_mioi
      (
      .this_val(accum_inter_0_5_val),
      .this_rdy(accum_inter_0_5_rdy),
      .this_msg(accum_inter_0_5_msg),
      .return_rsc_z(accum_inter_PushNB_5_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_6_mioi
      (
      .this_val(accum_inter_0_6_val),
      .this_rdy(accum_inter_0_6_rdy),
      .this_msg(accum_inter_0_6_msg),
      .return_rsc_z(accum_inter_PushNB_6_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  Connections_Combinational_SysPE_AccumType_Connections_SYN_PORT_PushNB  accum_inter_PushNB_7_mioi
      (
      .this_val(accum_inter_0_7_val),
      .this_rdy(accum_inter_0_7_rdy),
      .this_msg(accum_inter_0_7_msg),
      .return_rsc_z(accum_inter_PushNB_7_mioi_return_rsc_z),
      .ccs_MIO_clk(clk),
      .ccs_MIO_arst(rst),
      .ccs_ccore_start_rsc_dat(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  SysPE SysPE_1 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_0_val),
      .weight_in_rdy(weight_in_vec_0_rdy),
      .weight_in_msg(weight_in_vec_0_msg),
      .act_in_val(act_in_vec_0_val),
      .act_in_rdy(act_in_vec_0_rdy),
      .act_in_msg(act_in_vec_0_msg),
      .accum_in_val(accum_inter_0_0_val),
      .accum_in_rdy(accum_inter_0_0_rdy),
      .accum_in_msg(accum_inter_0_0_msg),
      .act_out_val(act_inter_0_0_val),
      .act_out_rdy(act_inter_0_0_rdy),
      .act_out_msg(act_inter_0_0_msg),
      .accum_out_val(accum_inter_1_0_val),
      .accum_out_rdy(accum_inter_1_0_rdy),
      .accum_out_msg(accum_inter_1_0_msg),
      .weight_out_val(weight_inter_0_0_val),
      .weight_out_rdy(weight_inter_0_0_rdy),
      .weight_out_msg(weight_inter_0_0_msg)
    );
  SysPE SysPE_1_1 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_1_val),
      .weight_in_rdy(weight_in_vec_1_rdy),
      .weight_in_msg(weight_in_vec_1_msg),
      .act_in_val(act_inter_0_0_val),
      .act_in_rdy(act_inter_0_0_rdy),
      .act_in_msg(act_inter_0_0_msg),
      .accum_in_val(accum_inter_0_1_val),
      .accum_in_rdy(accum_inter_0_1_rdy),
      .accum_in_msg(accum_inter_0_1_msg),
      .act_out_val(act_inter_0_1_val),
      .act_out_rdy(act_inter_0_1_rdy),
      .act_out_msg(act_inter_0_1_msg),
      .accum_out_val(accum_inter_1_1_val),
      .accum_out_rdy(accum_inter_1_1_rdy),
      .accum_out_msg(accum_inter_1_1_msg),
      .weight_out_val(weight_inter_0_1_val),
      .weight_out_rdy(weight_inter_0_1_rdy),
      .weight_out_msg(weight_inter_0_1_msg)
    );
  SysPE SysPE_2 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_2_val),
      .weight_in_rdy(weight_in_vec_2_rdy),
      .weight_in_msg(weight_in_vec_2_msg),
      .act_in_val(act_inter_0_1_val),
      .act_in_rdy(act_inter_0_1_rdy),
      .act_in_msg(act_inter_0_1_msg),
      .accum_in_val(accum_inter_0_2_val),
      .accum_in_rdy(accum_inter_0_2_rdy),
      .accum_in_msg(accum_inter_0_2_msg),
      .act_out_val(act_inter_0_2_val),
      .act_out_rdy(act_inter_0_2_rdy),
      .act_out_msg(act_inter_0_2_msg),
      .accum_out_val(accum_inter_1_2_val),
      .accum_out_rdy(accum_inter_1_2_rdy),
      .accum_out_msg(accum_inter_1_2_msg),
      .weight_out_val(weight_inter_0_2_val),
      .weight_out_rdy(weight_inter_0_2_rdy),
      .weight_out_msg(weight_inter_0_2_msg)
    );
  SysPE SysPE_3 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_3_val),
      .weight_in_rdy(weight_in_vec_3_rdy),
      .weight_in_msg(weight_in_vec_3_msg),
      .act_in_val(act_inter_0_2_val),
      .act_in_rdy(act_inter_0_2_rdy),
      .act_in_msg(act_inter_0_2_msg),
      .accum_in_val(accum_inter_0_3_val),
      .accum_in_rdy(accum_inter_0_3_rdy),
      .accum_in_msg(accum_inter_0_3_msg),
      .act_out_val(act_inter_0_3_val),
      .act_out_rdy(act_inter_0_3_rdy),
      .act_out_msg(act_inter_0_3_msg),
      .accum_out_val(accum_inter_1_3_val),
      .accum_out_rdy(accum_inter_1_3_rdy),
      .accum_out_msg(accum_inter_1_3_msg),
      .weight_out_val(weight_inter_0_3_val),
      .weight_out_rdy(weight_inter_0_3_rdy),
      .weight_out_msg(weight_inter_0_3_msg)
    );
  SysPE SysPE_4 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_4_val),
      .weight_in_rdy(weight_in_vec_4_rdy),
      .weight_in_msg(weight_in_vec_4_msg),
      .act_in_val(act_inter_0_3_val),
      .act_in_rdy(act_inter_0_3_rdy),
      .act_in_msg(act_inter_0_3_msg),
      .accum_in_val(accum_inter_0_4_val),
      .accum_in_rdy(accum_inter_0_4_rdy),
      .accum_in_msg(accum_inter_0_4_msg),
      .act_out_val(act_inter_0_4_val),
      .act_out_rdy(act_inter_0_4_rdy),
      .act_out_msg(act_inter_0_4_msg),
      .accum_out_val(accum_inter_1_4_val),
      .accum_out_rdy(accum_inter_1_4_rdy),
      .accum_out_msg(accum_inter_1_4_msg),
      .weight_out_val(weight_inter_0_4_val),
      .weight_out_rdy(weight_inter_0_4_rdy),
      .weight_out_msg(weight_inter_0_4_msg)
    );
  SysPE SysPE_5 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_5_val),
      .weight_in_rdy(weight_in_vec_5_rdy),
      .weight_in_msg(weight_in_vec_5_msg),
      .act_in_val(act_inter_0_4_val),
      .act_in_rdy(act_inter_0_4_rdy),
      .act_in_msg(act_inter_0_4_msg),
      .accum_in_val(accum_inter_0_5_val),
      .accum_in_rdy(accum_inter_0_5_rdy),
      .accum_in_msg(accum_inter_0_5_msg),
      .act_out_val(act_inter_0_5_val),
      .act_out_rdy(act_inter_0_5_rdy),
      .act_out_msg(act_inter_0_5_msg),
      .accum_out_val(accum_inter_1_5_val),
      .accum_out_rdy(accum_inter_1_5_rdy),
      .accum_out_msg(accum_inter_1_5_msg),
      .weight_out_val(weight_inter_0_5_val),
      .weight_out_rdy(weight_inter_0_5_rdy),
      .weight_out_msg(weight_inter_0_5_msg)
    );
  SysPE SysPE_6 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_6_val),
      .weight_in_rdy(weight_in_vec_6_rdy),
      .weight_in_msg(weight_in_vec_6_msg),
      .act_in_val(act_inter_0_5_val),
      .act_in_rdy(act_inter_0_5_rdy),
      .act_in_msg(act_inter_0_5_msg),
      .accum_in_val(accum_inter_0_6_val),
      .accum_in_rdy(accum_inter_0_6_rdy),
      .accum_in_msg(accum_inter_0_6_msg),
      .act_out_val(act_inter_0_6_val),
      .act_out_rdy(act_inter_0_6_rdy),
      .act_out_msg(act_inter_0_6_msg),
      .accum_out_val(accum_inter_1_6_val),
      .accum_out_rdy(accum_inter_1_6_rdy),
      .accum_out_msg(accum_inter_1_6_msg),
      .weight_out_val(weight_inter_0_6_val),
      .weight_out_rdy(weight_inter_0_6_rdy),
      .weight_out_msg(weight_inter_0_6_msg)
    );
  SysPE SysPE_7 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_in_vec_7_val),
      .weight_in_rdy(weight_in_vec_7_rdy),
      .weight_in_msg(weight_in_vec_7_msg),
      .act_in_val(act_inter_0_6_val),
      .act_in_rdy(act_inter_0_6_rdy),
      .act_in_msg(act_inter_0_6_msg),
      .accum_in_val(accum_inter_0_7_val),
      .accum_in_rdy(accum_inter_0_7_rdy),
      .accum_in_msg(accum_inter_0_7_msg),
      .act_out_val(act_inter_0_7_val),
      .act_out_rdy(act_inter_0_7_rdy),
      .act_out_msg(act_inter_0_7_msg),
      .accum_out_val(accum_inter_1_7_val),
      .accum_out_rdy(accum_inter_1_7_rdy),
      .accum_out_msg(accum_inter_1_7_msg),
      .weight_out_val(weight_inter_0_7_val),
      .weight_out_rdy(weight_inter_0_7_rdy),
      .weight_out_msg(weight_inter_0_7_msg)
    );
  SysPE SysPE_8 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_0_val),
      .weight_in_rdy(weight_inter_0_0_rdy),
      .weight_in_msg(weight_inter_0_0_msg),
      .act_in_val(act_in_vec_1_val),
      .act_in_rdy(act_in_vec_1_rdy),
      .act_in_msg(act_in_vec_1_msg),
      .accum_in_val(accum_inter_1_0_val),
      .accum_in_rdy(accum_inter_1_0_rdy),
      .accum_in_msg(accum_inter_1_0_msg),
      .act_out_val(act_inter_1_0_val),
      .act_out_rdy(act_inter_1_0_rdy),
      .act_out_msg(act_inter_1_0_msg),
      .accum_out_val(accum_inter_2_0_val),
      .accum_out_rdy(accum_inter_2_0_rdy),
      .accum_out_msg(accum_inter_2_0_msg),
      .weight_out_val(weight_inter_1_0_val),
      .weight_out_rdy(weight_inter_1_0_rdy),
      .weight_out_msg(weight_inter_1_0_msg)
    );
  SysPE SysPE_9 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_1_val),
      .weight_in_rdy(weight_inter_0_1_rdy),
      .weight_in_msg(weight_inter_0_1_msg),
      .act_in_val(act_inter_1_0_val),
      .act_in_rdy(act_inter_1_0_rdy),
      .act_in_msg(act_inter_1_0_msg),
      .accum_in_val(accum_inter_1_1_val),
      .accum_in_rdy(accum_inter_1_1_rdy),
      .accum_in_msg(accum_inter_1_1_msg),
      .act_out_val(act_inter_1_1_val),
      .act_out_rdy(act_inter_1_1_rdy),
      .act_out_msg(act_inter_1_1_msg),
      .accum_out_val(accum_inter_2_1_val),
      .accum_out_rdy(accum_inter_2_1_rdy),
      .accum_out_msg(accum_inter_2_1_msg),
      .weight_out_val(weight_inter_1_1_val),
      .weight_out_rdy(weight_inter_1_1_rdy),
      .weight_out_msg(weight_inter_1_1_msg)
    );
  SysPE SysPE_10 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_2_val),
      .weight_in_rdy(weight_inter_0_2_rdy),
      .weight_in_msg(weight_inter_0_2_msg),
      .act_in_val(act_inter_1_1_val),
      .act_in_rdy(act_inter_1_1_rdy),
      .act_in_msg(act_inter_1_1_msg),
      .accum_in_val(accum_inter_1_2_val),
      .accum_in_rdy(accum_inter_1_2_rdy),
      .accum_in_msg(accum_inter_1_2_msg),
      .act_out_val(act_inter_1_2_val),
      .act_out_rdy(act_inter_1_2_rdy),
      .act_out_msg(act_inter_1_2_msg),
      .accum_out_val(accum_inter_2_2_val),
      .accum_out_rdy(accum_inter_2_2_rdy),
      .accum_out_msg(accum_inter_2_2_msg),
      .weight_out_val(weight_inter_1_2_val),
      .weight_out_rdy(weight_inter_1_2_rdy),
      .weight_out_msg(weight_inter_1_2_msg)
    );
  SysPE SysPE_11 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_3_val),
      .weight_in_rdy(weight_inter_0_3_rdy),
      .weight_in_msg(weight_inter_0_3_msg),
      .act_in_val(act_inter_1_2_val),
      .act_in_rdy(act_inter_1_2_rdy),
      .act_in_msg(act_inter_1_2_msg),
      .accum_in_val(accum_inter_1_3_val),
      .accum_in_rdy(accum_inter_1_3_rdy),
      .accum_in_msg(accum_inter_1_3_msg),
      .act_out_val(act_inter_1_3_val),
      .act_out_rdy(act_inter_1_3_rdy),
      .act_out_msg(act_inter_1_3_msg),
      .accum_out_val(accum_inter_2_3_val),
      .accum_out_rdy(accum_inter_2_3_rdy),
      .accum_out_msg(accum_inter_2_3_msg),
      .weight_out_val(weight_inter_1_3_val),
      .weight_out_rdy(weight_inter_1_3_rdy),
      .weight_out_msg(weight_inter_1_3_msg)
    );
  SysPE SysPE_12 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_4_val),
      .weight_in_rdy(weight_inter_0_4_rdy),
      .weight_in_msg(weight_inter_0_4_msg),
      .act_in_val(act_inter_1_3_val),
      .act_in_rdy(act_inter_1_3_rdy),
      .act_in_msg(act_inter_1_3_msg),
      .accum_in_val(accum_inter_1_4_val),
      .accum_in_rdy(accum_inter_1_4_rdy),
      .accum_in_msg(accum_inter_1_4_msg),
      .act_out_val(act_inter_1_4_val),
      .act_out_rdy(act_inter_1_4_rdy),
      .act_out_msg(act_inter_1_4_msg),
      .accum_out_val(accum_inter_2_4_val),
      .accum_out_rdy(accum_inter_2_4_rdy),
      .accum_out_msg(accum_inter_2_4_msg),
      .weight_out_val(weight_inter_1_4_val),
      .weight_out_rdy(weight_inter_1_4_rdy),
      .weight_out_msg(weight_inter_1_4_msg)
    );
  SysPE SysPE_13 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_5_val),
      .weight_in_rdy(weight_inter_0_5_rdy),
      .weight_in_msg(weight_inter_0_5_msg),
      .act_in_val(act_inter_1_4_val),
      .act_in_rdy(act_inter_1_4_rdy),
      .act_in_msg(act_inter_1_4_msg),
      .accum_in_val(accum_inter_1_5_val),
      .accum_in_rdy(accum_inter_1_5_rdy),
      .accum_in_msg(accum_inter_1_5_msg),
      .act_out_val(act_inter_1_5_val),
      .act_out_rdy(act_inter_1_5_rdy),
      .act_out_msg(act_inter_1_5_msg),
      .accum_out_val(accum_inter_2_5_val),
      .accum_out_rdy(accum_inter_2_5_rdy),
      .accum_out_msg(accum_inter_2_5_msg),
      .weight_out_val(weight_inter_1_5_val),
      .weight_out_rdy(weight_inter_1_5_rdy),
      .weight_out_msg(weight_inter_1_5_msg)
    );
  SysPE SysPE_14 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_6_val),
      .weight_in_rdy(weight_inter_0_6_rdy),
      .weight_in_msg(weight_inter_0_6_msg),
      .act_in_val(act_inter_1_5_val),
      .act_in_rdy(act_inter_1_5_rdy),
      .act_in_msg(act_inter_1_5_msg),
      .accum_in_val(accum_inter_1_6_val),
      .accum_in_rdy(accum_inter_1_6_rdy),
      .accum_in_msg(accum_inter_1_6_msg),
      .act_out_val(act_inter_1_6_val),
      .act_out_rdy(act_inter_1_6_rdy),
      .act_out_msg(act_inter_1_6_msg),
      .accum_out_val(accum_inter_2_6_val),
      .accum_out_rdy(accum_inter_2_6_rdy),
      .accum_out_msg(accum_inter_2_6_msg),
      .weight_out_val(weight_inter_1_6_val),
      .weight_out_rdy(weight_inter_1_6_rdy),
      .weight_out_msg(weight_inter_1_6_msg)
    );
  SysPE SysPE_15 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_0_7_val),
      .weight_in_rdy(weight_inter_0_7_rdy),
      .weight_in_msg(weight_inter_0_7_msg),
      .act_in_val(act_inter_1_6_val),
      .act_in_rdy(act_inter_1_6_rdy),
      .act_in_msg(act_inter_1_6_msg),
      .accum_in_val(accum_inter_1_7_val),
      .accum_in_rdy(accum_inter_1_7_rdy),
      .accum_in_msg(accum_inter_1_7_msg),
      .act_out_val(act_inter_1_7_val),
      .act_out_rdy(act_inter_1_7_rdy),
      .act_out_msg(act_inter_1_7_msg),
      .accum_out_val(accum_inter_2_7_val),
      .accum_out_rdy(accum_inter_2_7_rdy),
      .accum_out_msg(accum_inter_2_7_msg),
      .weight_out_val(weight_inter_1_7_val),
      .weight_out_rdy(weight_inter_1_7_rdy),
      .weight_out_msg(weight_inter_1_7_msg)
    );
  SysPE SysPE_16 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_0_val),
      .weight_in_rdy(weight_inter_1_0_rdy),
      .weight_in_msg(weight_inter_1_0_msg),
      .act_in_val(act_in_vec_2_val),
      .act_in_rdy(act_in_vec_2_rdy),
      .act_in_msg(act_in_vec_2_msg),
      .accum_in_val(accum_inter_2_0_val),
      .accum_in_rdy(accum_inter_2_0_rdy),
      .accum_in_msg(accum_inter_2_0_msg),
      .act_out_val(act_inter_2_0_val),
      .act_out_rdy(act_inter_2_0_rdy),
      .act_out_msg(act_inter_2_0_msg),
      .accum_out_val(accum_inter_3_0_val),
      .accum_out_rdy(accum_inter_3_0_rdy),
      .accum_out_msg(accum_inter_3_0_msg),
      .weight_out_val(weight_inter_2_0_val),
      .weight_out_rdy(weight_inter_2_0_rdy),
      .weight_out_msg(weight_inter_2_0_msg)
    );
  SysPE SysPE_17 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_1_val),
      .weight_in_rdy(weight_inter_1_1_rdy),
      .weight_in_msg(weight_inter_1_1_msg),
      .act_in_val(act_inter_2_0_val),
      .act_in_rdy(act_inter_2_0_rdy),
      .act_in_msg(act_inter_2_0_msg),
      .accum_in_val(accum_inter_2_1_val),
      .accum_in_rdy(accum_inter_2_1_rdy),
      .accum_in_msg(accum_inter_2_1_msg),
      .act_out_val(act_inter_2_1_val),
      .act_out_rdy(act_inter_2_1_rdy),
      .act_out_msg(act_inter_2_1_msg),
      .accum_out_val(accum_inter_3_1_val),
      .accum_out_rdy(accum_inter_3_1_rdy),
      .accum_out_msg(accum_inter_3_1_msg),
      .weight_out_val(weight_inter_2_1_val),
      .weight_out_rdy(weight_inter_2_1_rdy),
      .weight_out_msg(weight_inter_2_1_msg)
    );
  SysPE SysPE_18 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_2_val),
      .weight_in_rdy(weight_inter_1_2_rdy),
      .weight_in_msg(weight_inter_1_2_msg),
      .act_in_val(act_inter_2_1_val),
      .act_in_rdy(act_inter_2_1_rdy),
      .act_in_msg(act_inter_2_1_msg),
      .accum_in_val(accum_inter_2_2_val),
      .accum_in_rdy(accum_inter_2_2_rdy),
      .accum_in_msg(accum_inter_2_2_msg),
      .act_out_val(act_inter_2_2_val),
      .act_out_rdy(act_inter_2_2_rdy),
      .act_out_msg(act_inter_2_2_msg),
      .accum_out_val(accum_inter_3_2_val),
      .accum_out_rdy(accum_inter_3_2_rdy),
      .accum_out_msg(accum_inter_3_2_msg),
      .weight_out_val(weight_inter_2_2_val),
      .weight_out_rdy(weight_inter_2_2_rdy),
      .weight_out_msg(weight_inter_2_2_msg)
    );
  SysPE SysPE_19 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_3_val),
      .weight_in_rdy(weight_inter_1_3_rdy),
      .weight_in_msg(weight_inter_1_3_msg),
      .act_in_val(act_inter_2_2_val),
      .act_in_rdy(act_inter_2_2_rdy),
      .act_in_msg(act_inter_2_2_msg),
      .accum_in_val(accum_inter_2_3_val),
      .accum_in_rdy(accum_inter_2_3_rdy),
      .accum_in_msg(accum_inter_2_3_msg),
      .act_out_val(act_inter_2_3_val),
      .act_out_rdy(act_inter_2_3_rdy),
      .act_out_msg(act_inter_2_3_msg),
      .accum_out_val(accum_inter_3_3_val),
      .accum_out_rdy(accum_inter_3_3_rdy),
      .accum_out_msg(accum_inter_3_3_msg),
      .weight_out_val(weight_inter_2_3_val),
      .weight_out_rdy(weight_inter_2_3_rdy),
      .weight_out_msg(weight_inter_2_3_msg)
    );
  SysPE SysPE_20 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_4_val),
      .weight_in_rdy(weight_inter_1_4_rdy),
      .weight_in_msg(weight_inter_1_4_msg),
      .act_in_val(act_inter_2_3_val),
      .act_in_rdy(act_inter_2_3_rdy),
      .act_in_msg(act_inter_2_3_msg),
      .accum_in_val(accum_inter_2_4_val),
      .accum_in_rdy(accum_inter_2_4_rdy),
      .accum_in_msg(accum_inter_2_4_msg),
      .act_out_val(act_inter_2_4_val),
      .act_out_rdy(act_inter_2_4_rdy),
      .act_out_msg(act_inter_2_4_msg),
      .accum_out_val(accum_inter_3_4_val),
      .accum_out_rdy(accum_inter_3_4_rdy),
      .accum_out_msg(accum_inter_3_4_msg),
      .weight_out_val(weight_inter_2_4_val),
      .weight_out_rdy(weight_inter_2_4_rdy),
      .weight_out_msg(weight_inter_2_4_msg)
    );
  SysPE SysPE_21 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_5_val),
      .weight_in_rdy(weight_inter_1_5_rdy),
      .weight_in_msg(weight_inter_1_5_msg),
      .act_in_val(act_inter_2_4_val),
      .act_in_rdy(act_inter_2_4_rdy),
      .act_in_msg(act_inter_2_4_msg),
      .accum_in_val(accum_inter_2_5_val),
      .accum_in_rdy(accum_inter_2_5_rdy),
      .accum_in_msg(accum_inter_2_5_msg),
      .act_out_val(act_inter_2_5_val),
      .act_out_rdy(act_inter_2_5_rdy),
      .act_out_msg(act_inter_2_5_msg),
      .accum_out_val(accum_inter_3_5_val),
      .accum_out_rdy(accum_inter_3_5_rdy),
      .accum_out_msg(accum_inter_3_5_msg),
      .weight_out_val(weight_inter_2_5_val),
      .weight_out_rdy(weight_inter_2_5_rdy),
      .weight_out_msg(weight_inter_2_5_msg)
    );
  SysPE SysPE_22 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_6_val),
      .weight_in_rdy(weight_inter_1_6_rdy),
      .weight_in_msg(weight_inter_1_6_msg),
      .act_in_val(act_inter_2_5_val),
      .act_in_rdy(act_inter_2_5_rdy),
      .act_in_msg(act_inter_2_5_msg),
      .accum_in_val(accum_inter_2_6_val),
      .accum_in_rdy(accum_inter_2_6_rdy),
      .accum_in_msg(accum_inter_2_6_msg),
      .act_out_val(act_inter_2_6_val),
      .act_out_rdy(act_inter_2_6_rdy),
      .act_out_msg(act_inter_2_6_msg),
      .accum_out_val(accum_inter_3_6_val),
      .accum_out_rdy(accum_inter_3_6_rdy),
      .accum_out_msg(accum_inter_3_6_msg),
      .weight_out_val(weight_inter_2_6_val),
      .weight_out_rdy(weight_inter_2_6_rdy),
      .weight_out_msg(weight_inter_2_6_msg)
    );
  SysPE SysPE_23 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_1_7_val),
      .weight_in_rdy(weight_inter_1_7_rdy),
      .weight_in_msg(weight_inter_1_7_msg),
      .act_in_val(act_inter_2_6_val),
      .act_in_rdy(act_inter_2_6_rdy),
      .act_in_msg(act_inter_2_6_msg),
      .accum_in_val(accum_inter_2_7_val),
      .accum_in_rdy(accum_inter_2_7_rdy),
      .accum_in_msg(accum_inter_2_7_msg),
      .act_out_val(act_inter_2_7_val),
      .act_out_rdy(act_inter_2_7_rdy),
      .act_out_msg(act_inter_2_7_msg),
      .accum_out_val(accum_inter_3_7_val),
      .accum_out_rdy(accum_inter_3_7_rdy),
      .accum_out_msg(accum_inter_3_7_msg),
      .weight_out_val(weight_inter_2_7_val),
      .weight_out_rdy(weight_inter_2_7_rdy),
      .weight_out_msg(weight_inter_2_7_msg)
    );
  SysPE SysPE_24 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_0_val),
      .weight_in_rdy(weight_inter_2_0_rdy),
      .weight_in_msg(weight_inter_2_0_msg),
      .act_in_val(act_in_vec_3_val),
      .act_in_rdy(act_in_vec_3_rdy),
      .act_in_msg(act_in_vec_3_msg),
      .accum_in_val(accum_inter_3_0_val),
      .accum_in_rdy(accum_inter_3_0_rdy),
      .accum_in_msg(accum_inter_3_0_msg),
      .act_out_val(act_inter_3_0_val),
      .act_out_rdy(act_inter_3_0_rdy),
      .act_out_msg(act_inter_3_0_msg),
      .accum_out_val(accum_inter_4_0_val),
      .accum_out_rdy(accum_inter_4_0_rdy),
      .accum_out_msg(accum_inter_4_0_msg),
      .weight_out_val(weight_inter_3_0_val),
      .weight_out_rdy(weight_inter_3_0_rdy),
      .weight_out_msg(weight_inter_3_0_msg)
    );
  SysPE SysPE_25 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_1_val),
      .weight_in_rdy(weight_inter_2_1_rdy),
      .weight_in_msg(weight_inter_2_1_msg),
      .act_in_val(act_inter_3_0_val),
      .act_in_rdy(act_inter_3_0_rdy),
      .act_in_msg(act_inter_3_0_msg),
      .accum_in_val(accum_inter_3_1_val),
      .accum_in_rdy(accum_inter_3_1_rdy),
      .accum_in_msg(accum_inter_3_1_msg),
      .act_out_val(act_inter_3_1_val),
      .act_out_rdy(act_inter_3_1_rdy),
      .act_out_msg(act_inter_3_1_msg),
      .accum_out_val(accum_inter_4_1_val),
      .accum_out_rdy(accum_inter_4_1_rdy),
      .accum_out_msg(accum_inter_4_1_msg),
      .weight_out_val(weight_inter_3_1_val),
      .weight_out_rdy(weight_inter_3_1_rdy),
      .weight_out_msg(weight_inter_3_1_msg)
    );
  SysPE SysPE_26 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_2_val),
      .weight_in_rdy(weight_inter_2_2_rdy),
      .weight_in_msg(weight_inter_2_2_msg),
      .act_in_val(act_inter_3_1_val),
      .act_in_rdy(act_inter_3_1_rdy),
      .act_in_msg(act_inter_3_1_msg),
      .accum_in_val(accum_inter_3_2_val),
      .accum_in_rdy(accum_inter_3_2_rdy),
      .accum_in_msg(accum_inter_3_2_msg),
      .act_out_val(act_inter_3_2_val),
      .act_out_rdy(act_inter_3_2_rdy),
      .act_out_msg(act_inter_3_2_msg),
      .accum_out_val(accum_inter_4_2_val),
      .accum_out_rdy(accum_inter_4_2_rdy),
      .accum_out_msg(accum_inter_4_2_msg),
      .weight_out_val(weight_inter_3_2_val),
      .weight_out_rdy(weight_inter_3_2_rdy),
      .weight_out_msg(weight_inter_3_2_msg)
    );
  SysPE SysPE_27 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_3_val),
      .weight_in_rdy(weight_inter_2_3_rdy),
      .weight_in_msg(weight_inter_2_3_msg),
      .act_in_val(act_inter_3_2_val),
      .act_in_rdy(act_inter_3_2_rdy),
      .act_in_msg(act_inter_3_2_msg),
      .accum_in_val(accum_inter_3_3_val),
      .accum_in_rdy(accum_inter_3_3_rdy),
      .accum_in_msg(accum_inter_3_3_msg),
      .act_out_val(act_inter_3_3_val),
      .act_out_rdy(act_inter_3_3_rdy),
      .act_out_msg(act_inter_3_3_msg),
      .accum_out_val(accum_inter_4_3_val),
      .accum_out_rdy(accum_inter_4_3_rdy),
      .accum_out_msg(accum_inter_4_3_msg),
      .weight_out_val(weight_inter_3_3_val),
      .weight_out_rdy(weight_inter_3_3_rdy),
      .weight_out_msg(weight_inter_3_3_msg)
    );
  SysPE SysPE_28 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_4_val),
      .weight_in_rdy(weight_inter_2_4_rdy),
      .weight_in_msg(weight_inter_2_4_msg),
      .act_in_val(act_inter_3_3_val),
      .act_in_rdy(act_inter_3_3_rdy),
      .act_in_msg(act_inter_3_3_msg),
      .accum_in_val(accum_inter_3_4_val),
      .accum_in_rdy(accum_inter_3_4_rdy),
      .accum_in_msg(accum_inter_3_4_msg),
      .act_out_val(act_inter_3_4_val),
      .act_out_rdy(act_inter_3_4_rdy),
      .act_out_msg(act_inter_3_4_msg),
      .accum_out_val(accum_inter_4_4_val),
      .accum_out_rdy(accum_inter_4_4_rdy),
      .accum_out_msg(accum_inter_4_4_msg),
      .weight_out_val(weight_inter_3_4_val),
      .weight_out_rdy(weight_inter_3_4_rdy),
      .weight_out_msg(weight_inter_3_4_msg)
    );
  SysPE SysPE_29 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_5_val),
      .weight_in_rdy(weight_inter_2_5_rdy),
      .weight_in_msg(weight_inter_2_5_msg),
      .act_in_val(act_inter_3_4_val),
      .act_in_rdy(act_inter_3_4_rdy),
      .act_in_msg(act_inter_3_4_msg),
      .accum_in_val(accum_inter_3_5_val),
      .accum_in_rdy(accum_inter_3_5_rdy),
      .accum_in_msg(accum_inter_3_5_msg),
      .act_out_val(act_inter_3_5_val),
      .act_out_rdy(act_inter_3_5_rdy),
      .act_out_msg(act_inter_3_5_msg),
      .accum_out_val(accum_inter_4_5_val),
      .accum_out_rdy(accum_inter_4_5_rdy),
      .accum_out_msg(accum_inter_4_5_msg),
      .weight_out_val(weight_inter_3_5_val),
      .weight_out_rdy(weight_inter_3_5_rdy),
      .weight_out_msg(weight_inter_3_5_msg)
    );
  SysPE SysPE_30 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_6_val),
      .weight_in_rdy(weight_inter_2_6_rdy),
      .weight_in_msg(weight_inter_2_6_msg),
      .act_in_val(act_inter_3_5_val),
      .act_in_rdy(act_inter_3_5_rdy),
      .act_in_msg(act_inter_3_5_msg),
      .accum_in_val(accum_inter_3_6_val),
      .accum_in_rdy(accum_inter_3_6_rdy),
      .accum_in_msg(accum_inter_3_6_msg),
      .act_out_val(act_inter_3_6_val),
      .act_out_rdy(act_inter_3_6_rdy),
      .act_out_msg(act_inter_3_6_msg),
      .accum_out_val(accum_inter_4_6_val),
      .accum_out_rdy(accum_inter_4_6_rdy),
      .accum_out_msg(accum_inter_4_6_msg),
      .weight_out_val(weight_inter_3_6_val),
      .weight_out_rdy(weight_inter_3_6_rdy),
      .weight_out_msg(weight_inter_3_6_msg)
    );
  SysPE SysPE_31 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_2_7_val),
      .weight_in_rdy(weight_inter_2_7_rdy),
      .weight_in_msg(weight_inter_2_7_msg),
      .act_in_val(act_inter_3_6_val),
      .act_in_rdy(act_inter_3_6_rdy),
      .act_in_msg(act_inter_3_6_msg),
      .accum_in_val(accum_inter_3_7_val),
      .accum_in_rdy(accum_inter_3_7_rdy),
      .accum_in_msg(accum_inter_3_7_msg),
      .act_out_val(act_inter_3_7_val),
      .act_out_rdy(act_inter_3_7_rdy),
      .act_out_msg(act_inter_3_7_msg),
      .accum_out_val(accum_inter_4_7_val),
      .accum_out_rdy(accum_inter_4_7_rdy),
      .accum_out_msg(accum_inter_4_7_msg),
      .weight_out_val(weight_inter_3_7_val),
      .weight_out_rdy(weight_inter_3_7_rdy),
      .weight_out_msg(weight_inter_3_7_msg)
    );
  SysPE SysPE_32 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_0_val),
      .weight_in_rdy(weight_inter_3_0_rdy),
      .weight_in_msg(weight_inter_3_0_msg),
      .act_in_val(act_in_vec_4_val),
      .act_in_rdy(act_in_vec_4_rdy),
      .act_in_msg(act_in_vec_4_msg),
      .accum_in_val(accum_inter_4_0_val),
      .accum_in_rdy(accum_inter_4_0_rdy),
      .accum_in_msg(accum_inter_4_0_msg),
      .act_out_val(act_inter_4_0_val),
      .act_out_rdy(act_inter_4_0_rdy),
      .act_out_msg(act_inter_4_0_msg),
      .accum_out_val(accum_inter_5_0_val),
      .accum_out_rdy(accum_inter_5_0_rdy),
      .accum_out_msg(accum_inter_5_0_msg),
      .weight_out_val(weight_inter_4_0_val),
      .weight_out_rdy(weight_inter_4_0_rdy),
      .weight_out_msg(weight_inter_4_0_msg)
    );
  SysPE SysPE_33 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_1_val),
      .weight_in_rdy(weight_inter_3_1_rdy),
      .weight_in_msg(weight_inter_3_1_msg),
      .act_in_val(act_inter_4_0_val),
      .act_in_rdy(act_inter_4_0_rdy),
      .act_in_msg(act_inter_4_0_msg),
      .accum_in_val(accum_inter_4_1_val),
      .accum_in_rdy(accum_inter_4_1_rdy),
      .accum_in_msg(accum_inter_4_1_msg),
      .act_out_val(act_inter_4_1_val),
      .act_out_rdy(act_inter_4_1_rdy),
      .act_out_msg(act_inter_4_1_msg),
      .accum_out_val(accum_inter_5_1_val),
      .accum_out_rdy(accum_inter_5_1_rdy),
      .accum_out_msg(accum_inter_5_1_msg),
      .weight_out_val(weight_inter_4_1_val),
      .weight_out_rdy(weight_inter_4_1_rdy),
      .weight_out_msg(weight_inter_4_1_msg)
    );
  SysPE SysPE_34 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_2_val),
      .weight_in_rdy(weight_inter_3_2_rdy),
      .weight_in_msg(weight_inter_3_2_msg),
      .act_in_val(act_inter_4_1_val),
      .act_in_rdy(act_inter_4_1_rdy),
      .act_in_msg(act_inter_4_1_msg),
      .accum_in_val(accum_inter_4_2_val),
      .accum_in_rdy(accum_inter_4_2_rdy),
      .accum_in_msg(accum_inter_4_2_msg),
      .act_out_val(act_inter_4_2_val),
      .act_out_rdy(act_inter_4_2_rdy),
      .act_out_msg(act_inter_4_2_msg),
      .accum_out_val(accum_inter_5_2_val),
      .accum_out_rdy(accum_inter_5_2_rdy),
      .accum_out_msg(accum_inter_5_2_msg),
      .weight_out_val(weight_inter_4_2_val),
      .weight_out_rdy(weight_inter_4_2_rdy),
      .weight_out_msg(weight_inter_4_2_msg)
    );
  SysPE SysPE_35 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_3_val),
      .weight_in_rdy(weight_inter_3_3_rdy),
      .weight_in_msg(weight_inter_3_3_msg),
      .act_in_val(act_inter_4_2_val),
      .act_in_rdy(act_inter_4_2_rdy),
      .act_in_msg(act_inter_4_2_msg),
      .accum_in_val(accum_inter_4_3_val),
      .accum_in_rdy(accum_inter_4_3_rdy),
      .accum_in_msg(accum_inter_4_3_msg),
      .act_out_val(act_inter_4_3_val),
      .act_out_rdy(act_inter_4_3_rdy),
      .act_out_msg(act_inter_4_3_msg),
      .accum_out_val(accum_inter_5_3_val),
      .accum_out_rdy(accum_inter_5_3_rdy),
      .accum_out_msg(accum_inter_5_3_msg),
      .weight_out_val(weight_inter_4_3_val),
      .weight_out_rdy(weight_inter_4_3_rdy),
      .weight_out_msg(weight_inter_4_3_msg)
    );
  SysPE SysPE_36 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_4_val),
      .weight_in_rdy(weight_inter_3_4_rdy),
      .weight_in_msg(weight_inter_3_4_msg),
      .act_in_val(act_inter_4_3_val),
      .act_in_rdy(act_inter_4_3_rdy),
      .act_in_msg(act_inter_4_3_msg),
      .accum_in_val(accum_inter_4_4_val),
      .accum_in_rdy(accum_inter_4_4_rdy),
      .accum_in_msg(accum_inter_4_4_msg),
      .act_out_val(act_inter_4_4_val),
      .act_out_rdy(act_inter_4_4_rdy),
      .act_out_msg(act_inter_4_4_msg),
      .accum_out_val(accum_inter_5_4_val),
      .accum_out_rdy(accum_inter_5_4_rdy),
      .accum_out_msg(accum_inter_5_4_msg),
      .weight_out_val(weight_inter_4_4_val),
      .weight_out_rdy(weight_inter_4_4_rdy),
      .weight_out_msg(weight_inter_4_4_msg)
    );
  SysPE SysPE_37 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_5_val),
      .weight_in_rdy(weight_inter_3_5_rdy),
      .weight_in_msg(weight_inter_3_5_msg),
      .act_in_val(act_inter_4_4_val),
      .act_in_rdy(act_inter_4_4_rdy),
      .act_in_msg(act_inter_4_4_msg),
      .accum_in_val(accum_inter_4_5_val),
      .accum_in_rdy(accum_inter_4_5_rdy),
      .accum_in_msg(accum_inter_4_5_msg),
      .act_out_val(act_inter_4_5_val),
      .act_out_rdy(act_inter_4_5_rdy),
      .act_out_msg(act_inter_4_5_msg),
      .accum_out_val(accum_inter_5_5_val),
      .accum_out_rdy(accum_inter_5_5_rdy),
      .accum_out_msg(accum_inter_5_5_msg),
      .weight_out_val(weight_inter_4_5_val),
      .weight_out_rdy(weight_inter_4_5_rdy),
      .weight_out_msg(weight_inter_4_5_msg)
    );
  SysPE SysPE_38 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_6_val),
      .weight_in_rdy(weight_inter_3_6_rdy),
      .weight_in_msg(weight_inter_3_6_msg),
      .act_in_val(act_inter_4_5_val),
      .act_in_rdy(act_inter_4_5_rdy),
      .act_in_msg(act_inter_4_5_msg),
      .accum_in_val(accum_inter_4_6_val),
      .accum_in_rdy(accum_inter_4_6_rdy),
      .accum_in_msg(accum_inter_4_6_msg),
      .act_out_val(act_inter_4_6_val),
      .act_out_rdy(act_inter_4_6_rdy),
      .act_out_msg(act_inter_4_6_msg),
      .accum_out_val(accum_inter_5_6_val),
      .accum_out_rdy(accum_inter_5_6_rdy),
      .accum_out_msg(accum_inter_5_6_msg),
      .weight_out_val(weight_inter_4_6_val),
      .weight_out_rdy(weight_inter_4_6_rdy),
      .weight_out_msg(weight_inter_4_6_msg)
    );
  SysPE SysPE_39 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_3_7_val),
      .weight_in_rdy(weight_inter_3_7_rdy),
      .weight_in_msg(weight_inter_3_7_msg),
      .act_in_val(act_inter_4_6_val),
      .act_in_rdy(act_inter_4_6_rdy),
      .act_in_msg(act_inter_4_6_msg),
      .accum_in_val(accum_inter_4_7_val),
      .accum_in_rdy(accum_inter_4_7_rdy),
      .accum_in_msg(accum_inter_4_7_msg),
      .act_out_val(act_inter_4_7_val),
      .act_out_rdy(act_inter_4_7_rdy),
      .act_out_msg(act_inter_4_7_msg),
      .accum_out_val(accum_inter_5_7_val),
      .accum_out_rdy(accum_inter_5_7_rdy),
      .accum_out_msg(accum_inter_5_7_msg),
      .weight_out_val(weight_inter_4_7_val),
      .weight_out_rdy(weight_inter_4_7_rdy),
      .weight_out_msg(weight_inter_4_7_msg)
    );
  SysPE SysPE_40 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_0_val),
      .weight_in_rdy(weight_inter_4_0_rdy),
      .weight_in_msg(weight_inter_4_0_msg),
      .act_in_val(act_in_vec_5_val),
      .act_in_rdy(act_in_vec_5_rdy),
      .act_in_msg(act_in_vec_5_msg),
      .accum_in_val(accum_inter_5_0_val),
      .accum_in_rdy(accum_inter_5_0_rdy),
      .accum_in_msg(accum_inter_5_0_msg),
      .act_out_val(act_inter_5_0_val),
      .act_out_rdy(act_inter_5_0_rdy),
      .act_out_msg(act_inter_5_0_msg),
      .accum_out_val(accum_inter_6_0_val),
      .accum_out_rdy(accum_inter_6_0_rdy),
      .accum_out_msg(accum_inter_6_0_msg),
      .weight_out_val(weight_inter_5_0_val),
      .weight_out_rdy(weight_inter_5_0_rdy),
      .weight_out_msg(weight_inter_5_0_msg)
    );
  SysPE SysPE_41 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_1_val),
      .weight_in_rdy(weight_inter_4_1_rdy),
      .weight_in_msg(weight_inter_4_1_msg),
      .act_in_val(act_inter_5_0_val),
      .act_in_rdy(act_inter_5_0_rdy),
      .act_in_msg(act_inter_5_0_msg),
      .accum_in_val(accum_inter_5_1_val),
      .accum_in_rdy(accum_inter_5_1_rdy),
      .accum_in_msg(accum_inter_5_1_msg),
      .act_out_val(act_inter_5_1_val),
      .act_out_rdy(act_inter_5_1_rdy),
      .act_out_msg(act_inter_5_1_msg),
      .accum_out_val(accum_inter_6_1_val),
      .accum_out_rdy(accum_inter_6_1_rdy),
      .accum_out_msg(accum_inter_6_1_msg),
      .weight_out_val(weight_inter_5_1_val),
      .weight_out_rdy(weight_inter_5_1_rdy),
      .weight_out_msg(weight_inter_5_1_msg)
    );
  SysPE SysPE_42 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_2_val),
      .weight_in_rdy(weight_inter_4_2_rdy),
      .weight_in_msg(weight_inter_4_2_msg),
      .act_in_val(act_inter_5_1_val),
      .act_in_rdy(act_inter_5_1_rdy),
      .act_in_msg(act_inter_5_1_msg),
      .accum_in_val(accum_inter_5_2_val),
      .accum_in_rdy(accum_inter_5_2_rdy),
      .accum_in_msg(accum_inter_5_2_msg),
      .act_out_val(act_inter_5_2_val),
      .act_out_rdy(act_inter_5_2_rdy),
      .act_out_msg(act_inter_5_2_msg),
      .accum_out_val(accum_inter_6_2_val),
      .accum_out_rdy(accum_inter_6_2_rdy),
      .accum_out_msg(accum_inter_6_2_msg),
      .weight_out_val(weight_inter_5_2_val),
      .weight_out_rdy(weight_inter_5_2_rdy),
      .weight_out_msg(weight_inter_5_2_msg)
    );
  SysPE SysPE_43 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_3_val),
      .weight_in_rdy(weight_inter_4_3_rdy),
      .weight_in_msg(weight_inter_4_3_msg),
      .act_in_val(act_inter_5_2_val),
      .act_in_rdy(act_inter_5_2_rdy),
      .act_in_msg(act_inter_5_2_msg),
      .accum_in_val(accum_inter_5_3_val),
      .accum_in_rdy(accum_inter_5_3_rdy),
      .accum_in_msg(accum_inter_5_3_msg),
      .act_out_val(act_inter_5_3_val),
      .act_out_rdy(act_inter_5_3_rdy),
      .act_out_msg(act_inter_5_3_msg),
      .accum_out_val(accum_inter_6_3_val),
      .accum_out_rdy(accum_inter_6_3_rdy),
      .accum_out_msg(accum_inter_6_3_msg),
      .weight_out_val(weight_inter_5_3_val),
      .weight_out_rdy(weight_inter_5_3_rdy),
      .weight_out_msg(weight_inter_5_3_msg)
    );
  SysPE SysPE_44 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_4_val),
      .weight_in_rdy(weight_inter_4_4_rdy),
      .weight_in_msg(weight_inter_4_4_msg),
      .act_in_val(act_inter_5_3_val),
      .act_in_rdy(act_inter_5_3_rdy),
      .act_in_msg(act_inter_5_3_msg),
      .accum_in_val(accum_inter_5_4_val),
      .accum_in_rdy(accum_inter_5_4_rdy),
      .accum_in_msg(accum_inter_5_4_msg),
      .act_out_val(act_inter_5_4_val),
      .act_out_rdy(act_inter_5_4_rdy),
      .act_out_msg(act_inter_5_4_msg),
      .accum_out_val(accum_inter_6_4_val),
      .accum_out_rdy(accum_inter_6_4_rdy),
      .accum_out_msg(accum_inter_6_4_msg),
      .weight_out_val(weight_inter_5_4_val),
      .weight_out_rdy(weight_inter_5_4_rdy),
      .weight_out_msg(weight_inter_5_4_msg)
    );
  SysPE SysPE_45 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_5_val),
      .weight_in_rdy(weight_inter_4_5_rdy),
      .weight_in_msg(weight_inter_4_5_msg),
      .act_in_val(act_inter_5_4_val),
      .act_in_rdy(act_inter_5_4_rdy),
      .act_in_msg(act_inter_5_4_msg),
      .accum_in_val(accum_inter_5_5_val),
      .accum_in_rdy(accum_inter_5_5_rdy),
      .accum_in_msg(accum_inter_5_5_msg),
      .act_out_val(act_inter_5_5_val),
      .act_out_rdy(act_inter_5_5_rdy),
      .act_out_msg(act_inter_5_5_msg),
      .accum_out_val(accum_inter_6_5_val),
      .accum_out_rdy(accum_inter_6_5_rdy),
      .accum_out_msg(accum_inter_6_5_msg),
      .weight_out_val(weight_inter_5_5_val),
      .weight_out_rdy(weight_inter_5_5_rdy),
      .weight_out_msg(weight_inter_5_5_msg)
    );
  SysPE SysPE_46 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_6_val),
      .weight_in_rdy(weight_inter_4_6_rdy),
      .weight_in_msg(weight_inter_4_6_msg),
      .act_in_val(act_inter_5_5_val),
      .act_in_rdy(act_inter_5_5_rdy),
      .act_in_msg(act_inter_5_5_msg),
      .accum_in_val(accum_inter_5_6_val),
      .accum_in_rdy(accum_inter_5_6_rdy),
      .accum_in_msg(accum_inter_5_6_msg),
      .act_out_val(act_inter_5_6_val),
      .act_out_rdy(act_inter_5_6_rdy),
      .act_out_msg(act_inter_5_6_msg),
      .accum_out_val(accum_inter_6_6_val),
      .accum_out_rdy(accum_inter_6_6_rdy),
      .accum_out_msg(accum_inter_6_6_msg),
      .weight_out_val(weight_inter_5_6_val),
      .weight_out_rdy(weight_inter_5_6_rdy),
      .weight_out_msg(weight_inter_5_6_msg)
    );
  SysPE SysPE_47 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_4_7_val),
      .weight_in_rdy(weight_inter_4_7_rdy),
      .weight_in_msg(weight_inter_4_7_msg),
      .act_in_val(act_inter_5_6_val),
      .act_in_rdy(act_inter_5_6_rdy),
      .act_in_msg(act_inter_5_6_msg),
      .accum_in_val(accum_inter_5_7_val),
      .accum_in_rdy(accum_inter_5_7_rdy),
      .accum_in_msg(accum_inter_5_7_msg),
      .act_out_val(act_inter_5_7_val),
      .act_out_rdy(act_inter_5_7_rdy),
      .act_out_msg(act_inter_5_7_msg),
      .accum_out_val(accum_inter_6_7_val),
      .accum_out_rdy(accum_inter_6_7_rdy),
      .accum_out_msg(accum_inter_6_7_msg),
      .weight_out_val(weight_inter_5_7_val),
      .weight_out_rdy(weight_inter_5_7_rdy),
      .weight_out_msg(weight_inter_5_7_msg)
    );
  SysPE SysPE_48 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_0_val),
      .weight_in_rdy(weight_inter_5_0_rdy),
      .weight_in_msg(weight_inter_5_0_msg),
      .act_in_val(act_in_vec_6_val),
      .act_in_rdy(act_in_vec_6_rdy),
      .act_in_msg(act_in_vec_6_msg),
      .accum_in_val(accum_inter_6_0_val),
      .accum_in_rdy(accum_inter_6_0_rdy),
      .accum_in_msg(accum_inter_6_0_msg),
      .act_out_val(act_inter_6_0_val),
      .act_out_rdy(act_inter_6_0_rdy),
      .act_out_msg(act_inter_6_0_msg),
      .accum_out_val(accum_inter_7_0_val),
      .accum_out_rdy(accum_inter_7_0_rdy),
      .accum_out_msg(accum_inter_7_0_msg),
      .weight_out_val(weight_inter_6_0_val),
      .weight_out_rdy(weight_inter_6_0_rdy),
      .weight_out_msg(weight_inter_6_0_msg)
    );
  SysPE SysPE_49 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_1_val),
      .weight_in_rdy(weight_inter_5_1_rdy),
      .weight_in_msg(weight_inter_5_1_msg),
      .act_in_val(act_inter_6_0_val),
      .act_in_rdy(act_inter_6_0_rdy),
      .act_in_msg(act_inter_6_0_msg),
      .accum_in_val(accum_inter_6_1_val),
      .accum_in_rdy(accum_inter_6_1_rdy),
      .accum_in_msg(accum_inter_6_1_msg),
      .act_out_val(act_inter_6_1_val),
      .act_out_rdy(act_inter_6_1_rdy),
      .act_out_msg(act_inter_6_1_msg),
      .accum_out_val(accum_inter_7_1_val),
      .accum_out_rdy(accum_inter_7_1_rdy),
      .accum_out_msg(accum_inter_7_1_msg),
      .weight_out_val(weight_inter_6_1_val),
      .weight_out_rdy(weight_inter_6_1_rdy),
      .weight_out_msg(weight_inter_6_1_msg)
    );
  SysPE SysPE_50 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_2_val),
      .weight_in_rdy(weight_inter_5_2_rdy),
      .weight_in_msg(weight_inter_5_2_msg),
      .act_in_val(act_inter_6_1_val),
      .act_in_rdy(act_inter_6_1_rdy),
      .act_in_msg(act_inter_6_1_msg),
      .accum_in_val(accum_inter_6_2_val),
      .accum_in_rdy(accum_inter_6_2_rdy),
      .accum_in_msg(accum_inter_6_2_msg),
      .act_out_val(act_inter_6_2_val),
      .act_out_rdy(act_inter_6_2_rdy),
      .act_out_msg(act_inter_6_2_msg),
      .accum_out_val(accum_inter_7_2_val),
      .accum_out_rdy(accum_inter_7_2_rdy),
      .accum_out_msg(accum_inter_7_2_msg),
      .weight_out_val(weight_inter_6_2_val),
      .weight_out_rdy(weight_inter_6_2_rdy),
      .weight_out_msg(weight_inter_6_2_msg)
    );
  SysPE SysPE_51 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_3_val),
      .weight_in_rdy(weight_inter_5_3_rdy),
      .weight_in_msg(weight_inter_5_3_msg),
      .act_in_val(act_inter_6_2_val),
      .act_in_rdy(act_inter_6_2_rdy),
      .act_in_msg(act_inter_6_2_msg),
      .accum_in_val(accum_inter_6_3_val),
      .accum_in_rdy(accum_inter_6_3_rdy),
      .accum_in_msg(accum_inter_6_3_msg),
      .act_out_val(act_inter_6_3_val),
      .act_out_rdy(act_inter_6_3_rdy),
      .act_out_msg(act_inter_6_3_msg),
      .accum_out_val(accum_inter_7_3_val),
      .accum_out_rdy(accum_inter_7_3_rdy),
      .accum_out_msg(accum_inter_7_3_msg),
      .weight_out_val(weight_inter_6_3_val),
      .weight_out_rdy(weight_inter_6_3_rdy),
      .weight_out_msg(weight_inter_6_3_msg)
    );
  SysPE SysPE_52 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_4_val),
      .weight_in_rdy(weight_inter_5_4_rdy),
      .weight_in_msg(weight_inter_5_4_msg),
      .act_in_val(act_inter_6_3_val),
      .act_in_rdy(act_inter_6_3_rdy),
      .act_in_msg(act_inter_6_3_msg),
      .accum_in_val(accum_inter_6_4_val),
      .accum_in_rdy(accum_inter_6_4_rdy),
      .accum_in_msg(accum_inter_6_4_msg),
      .act_out_val(act_inter_6_4_val),
      .act_out_rdy(act_inter_6_4_rdy),
      .act_out_msg(act_inter_6_4_msg),
      .accum_out_val(accum_inter_7_4_val),
      .accum_out_rdy(accum_inter_7_4_rdy),
      .accum_out_msg(accum_inter_7_4_msg),
      .weight_out_val(weight_inter_6_4_val),
      .weight_out_rdy(weight_inter_6_4_rdy),
      .weight_out_msg(weight_inter_6_4_msg)
    );
  SysPE SysPE_53 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_5_val),
      .weight_in_rdy(weight_inter_5_5_rdy),
      .weight_in_msg(weight_inter_5_5_msg),
      .act_in_val(act_inter_6_4_val),
      .act_in_rdy(act_inter_6_4_rdy),
      .act_in_msg(act_inter_6_4_msg),
      .accum_in_val(accum_inter_6_5_val),
      .accum_in_rdy(accum_inter_6_5_rdy),
      .accum_in_msg(accum_inter_6_5_msg),
      .act_out_val(act_inter_6_5_val),
      .act_out_rdy(act_inter_6_5_rdy),
      .act_out_msg(act_inter_6_5_msg),
      .accum_out_val(accum_inter_7_5_val),
      .accum_out_rdy(accum_inter_7_5_rdy),
      .accum_out_msg(accum_inter_7_5_msg),
      .weight_out_val(weight_inter_6_5_val),
      .weight_out_rdy(weight_inter_6_5_rdy),
      .weight_out_msg(weight_inter_6_5_msg)
    );
  SysPE SysPE_54 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_6_val),
      .weight_in_rdy(weight_inter_5_6_rdy),
      .weight_in_msg(weight_inter_5_6_msg),
      .act_in_val(act_inter_6_5_val),
      .act_in_rdy(act_inter_6_5_rdy),
      .act_in_msg(act_inter_6_5_msg),
      .accum_in_val(accum_inter_6_6_val),
      .accum_in_rdy(accum_inter_6_6_rdy),
      .accum_in_msg(accum_inter_6_6_msg),
      .act_out_val(act_inter_6_6_val),
      .act_out_rdy(act_inter_6_6_rdy),
      .act_out_msg(act_inter_6_6_msg),
      .accum_out_val(accum_inter_7_6_val),
      .accum_out_rdy(accum_inter_7_6_rdy),
      .accum_out_msg(accum_inter_7_6_msg),
      .weight_out_val(weight_inter_6_6_val),
      .weight_out_rdy(weight_inter_6_6_rdy),
      .weight_out_msg(weight_inter_6_6_msg)
    );
  SysPE SysPE_55 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_5_7_val),
      .weight_in_rdy(weight_inter_5_7_rdy),
      .weight_in_msg(weight_inter_5_7_msg),
      .act_in_val(act_inter_6_6_val),
      .act_in_rdy(act_inter_6_6_rdy),
      .act_in_msg(act_inter_6_6_msg),
      .accum_in_val(accum_inter_6_7_val),
      .accum_in_rdy(accum_inter_6_7_rdy),
      .accum_in_msg(accum_inter_6_7_msg),
      .act_out_val(act_inter_6_7_val),
      .act_out_rdy(act_inter_6_7_rdy),
      .act_out_msg(act_inter_6_7_msg),
      .accum_out_val(accum_inter_7_7_val),
      .accum_out_rdy(accum_inter_7_7_rdy),
      .accum_out_msg(accum_inter_7_7_msg),
      .weight_out_val(weight_inter_6_7_val),
      .weight_out_rdy(weight_inter_6_7_rdy),
      .weight_out_msg(weight_inter_6_7_msg)
    );
  SysPE SysPE_56 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_0_val),
      .weight_in_rdy(weight_inter_6_0_rdy),
      .weight_in_msg(weight_inter_6_0_msg),
      .act_in_val(act_in_vec_7_val),
      .act_in_rdy(act_in_vec_7_rdy),
      .act_in_msg(act_in_vec_7_msg),
      .accum_in_val(accum_inter_7_0_val),
      .accum_in_rdy(accum_inter_7_0_rdy),
      .accum_in_msg(accum_inter_7_0_msg),
      .act_out_val(act_inter_7_0_val),
      .act_out_rdy(act_inter_7_0_rdy),
      .act_out_msg(act_inter_7_0_msg),
      .accum_out_val(accum_out_vec_0_val),
      .accum_out_rdy(accum_out_vec_0_rdy),
      .accum_out_msg(accum_out_vec_0_msg),
      .weight_out_val(weight_inter_7_0_val),
      .weight_out_rdy(weight_inter_7_0_rdy),
      .weight_out_msg(weight_inter_7_0_msg)
    );
  SysPE SysPE_57 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_1_val),
      .weight_in_rdy(weight_inter_6_1_rdy),
      .weight_in_msg(weight_inter_6_1_msg),
      .act_in_val(act_inter_7_0_val),
      .act_in_rdy(act_inter_7_0_rdy),
      .act_in_msg(act_inter_7_0_msg),
      .accum_in_val(accum_inter_7_1_val),
      .accum_in_rdy(accum_inter_7_1_rdy),
      .accum_in_msg(accum_inter_7_1_msg),
      .act_out_val(act_inter_7_1_val),
      .act_out_rdy(act_inter_7_1_rdy),
      .act_out_msg(act_inter_7_1_msg),
      .accum_out_val(accum_out_vec_1_val),
      .accum_out_rdy(accum_out_vec_1_rdy),
      .accum_out_msg(accum_out_vec_1_msg),
      .weight_out_val(weight_inter_7_1_val),
      .weight_out_rdy(weight_inter_7_1_rdy),
      .weight_out_msg(weight_inter_7_1_msg)
    );
  SysPE SysPE_58 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_2_val),
      .weight_in_rdy(weight_inter_6_2_rdy),
      .weight_in_msg(weight_inter_6_2_msg),
      .act_in_val(act_inter_7_1_val),
      .act_in_rdy(act_inter_7_1_rdy),
      .act_in_msg(act_inter_7_1_msg),
      .accum_in_val(accum_inter_7_2_val),
      .accum_in_rdy(accum_inter_7_2_rdy),
      .accum_in_msg(accum_inter_7_2_msg),
      .act_out_val(act_inter_7_2_val),
      .act_out_rdy(act_inter_7_2_rdy),
      .act_out_msg(act_inter_7_2_msg),
      .accum_out_val(accum_out_vec_2_val),
      .accum_out_rdy(accum_out_vec_2_rdy),
      .accum_out_msg(accum_out_vec_2_msg),
      .weight_out_val(weight_inter_7_2_val),
      .weight_out_rdy(weight_inter_7_2_rdy),
      .weight_out_msg(weight_inter_7_2_msg)
    );
  SysPE SysPE_59 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_3_val),
      .weight_in_rdy(weight_inter_6_3_rdy),
      .weight_in_msg(weight_inter_6_3_msg),
      .act_in_val(act_inter_7_2_val),
      .act_in_rdy(act_inter_7_2_rdy),
      .act_in_msg(act_inter_7_2_msg),
      .accum_in_val(accum_inter_7_3_val),
      .accum_in_rdy(accum_inter_7_3_rdy),
      .accum_in_msg(accum_inter_7_3_msg),
      .act_out_val(act_inter_7_3_val),
      .act_out_rdy(act_inter_7_3_rdy),
      .act_out_msg(act_inter_7_3_msg),
      .accum_out_val(accum_out_vec_3_val),
      .accum_out_rdy(accum_out_vec_3_rdy),
      .accum_out_msg(accum_out_vec_3_msg),
      .weight_out_val(weight_inter_7_3_val),
      .weight_out_rdy(weight_inter_7_3_rdy),
      .weight_out_msg(weight_inter_7_3_msg)
    );
  SysPE SysPE_60 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_4_val),
      .weight_in_rdy(weight_inter_6_4_rdy),
      .weight_in_msg(weight_inter_6_4_msg),
      .act_in_val(act_inter_7_3_val),
      .act_in_rdy(act_inter_7_3_rdy),
      .act_in_msg(act_inter_7_3_msg),
      .accum_in_val(accum_inter_7_4_val),
      .accum_in_rdy(accum_inter_7_4_rdy),
      .accum_in_msg(accum_inter_7_4_msg),
      .act_out_val(act_inter_7_4_val),
      .act_out_rdy(act_inter_7_4_rdy),
      .act_out_msg(act_inter_7_4_msg),
      .accum_out_val(accum_out_vec_4_val),
      .accum_out_rdy(accum_out_vec_4_rdy),
      .accum_out_msg(accum_out_vec_4_msg),
      .weight_out_val(weight_inter_7_4_val),
      .weight_out_rdy(weight_inter_7_4_rdy),
      .weight_out_msg(weight_inter_7_4_msg)
    );
  SysPE SysPE_61 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_5_val),
      .weight_in_rdy(weight_inter_6_5_rdy),
      .weight_in_msg(weight_inter_6_5_msg),
      .act_in_val(act_inter_7_4_val),
      .act_in_rdy(act_inter_7_4_rdy),
      .act_in_msg(act_inter_7_4_msg),
      .accum_in_val(accum_inter_7_5_val),
      .accum_in_rdy(accum_inter_7_5_rdy),
      .accum_in_msg(accum_inter_7_5_msg),
      .act_out_val(act_inter_7_5_val),
      .act_out_rdy(act_inter_7_5_rdy),
      .act_out_msg(act_inter_7_5_msg),
      .accum_out_val(accum_out_vec_5_val),
      .accum_out_rdy(accum_out_vec_5_rdy),
      .accum_out_msg(accum_out_vec_5_msg),
      .weight_out_val(weight_inter_7_5_val),
      .weight_out_rdy(weight_inter_7_5_rdy),
      .weight_out_msg(weight_inter_7_5_msg)
    );
  SysPE SysPE_62 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_6_val),
      .weight_in_rdy(weight_inter_6_6_rdy),
      .weight_in_msg(weight_inter_6_6_msg),
      .act_in_val(act_inter_7_5_val),
      .act_in_rdy(act_inter_7_5_rdy),
      .act_in_msg(act_inter_7_5_msg),
      .accum_in_val(accum_inter_7_6_val),
      .accum_in_rdy(accum_inter_7_6_rdy),
      .accum_in_msg(accum_inter_7_6_msg),
      .act_out_val(act_inter_7_6_val),
      .act_out_rdy(act_inter_7_6_rdy),
      .act_out_msg(act_inter_7_6_msg),
      .accum_out_val(accum_out_vec_6_val),
      .accum_out_rdy(accum_out_vec_6_rdy),
      .accum_out_msg(accum_out_vec_6_msg),
      .weight_out_val(weight_inter_7_6_val),
      .weight_out_rdy(weight_inter_7_6_rdy),
      .weight_out_msg(weight_inter_7_6_msg)
    );
  SysPE SysPE_63 (
      .clk(clk),
      .rst(rst),
      .weight_in_val(weight_inter_6_7_val),
      .weight_in_rdy(weight_inter_6_7_rdy),
      .weight_in_msg(weight_inter_6_7_msg),
      .act_in_val(act_inter_7_6_val),
      .act_in_rdy(act_inter_7_6_rdy),
      .act_in_msg(act_inter_7_6_msg),
      .accum_in_val(accum_inter_7_7_val),
      .accum_in_rdy(accum_inter_7_7_rdy),
      .accum_in_msg(accum_inter_7_7_msg),
      .act_out_val(act_inter_7_7_val),
      .act_out_rdy(act_inter_7_7_rdy),
      .act_out_msg(act_inter_7_7_msg),
      .accum_out_val(accum_out_vec_7_val),
      .accum_out_rdy(accum_out_vec_7_rdy),
      .accum_out_msg(accum_out_vec_7_msg),
      .weight_out_val(weight_inter_7_7_val),
      .weight_out_rdy(weight_inter_7_7_rdy),
      .weight_out_msg(weight_inter_7_7_msg)
    );
  SysArray_WeightOutRun SysArray_WeightOutRun_inst (
      .clk(clk),
      .rst(rst),
      .weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_pff(weight_inter_PopNB_56_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  SysArray_ActOutRun SysArray_ActOutRun_inst (
      .clk(clk),
      .rst(rst),
      .act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_pff(act_inter_PopNB_7_mioi_ccs_ccore_start_rsc_dat_iff)
    );
  SysArray_AccumInRun SysArray_AccumInRun_inst (
      .clk(clk),
      .rst(rst),
      .accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_pff(accum_inter_PushNB_mioi_ccs_ccore_start_rsc_dat_iff)
    );
endmodule

// ------------------------------------------------------------------
//  Design Unit:    SysTop_rtl
// ------------------------------------------------------------------


module SysTop_rtl (
  clk, rst, write_req_val, write_req_rdy, write_req_msg, start_val, start_rdy, start_msg,
      weight_in_vec_0_val, weight_in_vec_1_val, weight_in_vec_2_val, weight_in_vec_3_val,
      weight_in_vec_4_val, weight_in_vec_5_val, weight_in_vec_6_val, weight_in_vec_7_val,
      weight_in_vec_0_rdy, weight_in_vec_1_rdy, weight_in_vec_2_rdy, weight_in_vec_3_rdy,
      weight_in_vec_4_rdy, weight_in_vec_5_rdy, weight_in_vec_6_rdy, weight_in_vec_7_rdy,
      weight_in_vec_0_msg, weight_in_vec_1_msg, weight_in_vec_2_msg, weight_in_vec_3_msg,
      weight_in_vec_4_msg, weight_in_vec_5_msg, weight_in_vec_6_msg, weight_in_vec_7_msg,
      accum_out_vec_0_val, accum_out_vec_1_val, accum_out_vec_2_val, accum_out_vec_3_val,
      accum_out_vec_4_val, accum_out_vec_5_val, accum_out_vec_6_val, accum_out_vec_7_val,
      accum_out_vec_0_rdy, accum_out_vec_1_rdy, accum_out_vec_2_rdy, accum_out_vec_3_rdy,
      accum_out_vec_4_rdy, accum_out_vec_5_rdy, accum_out_vec_6_rdy, accum_out_vec_7_rdy,
      accum_out_vec_0_msg, accum_out_vec_1_msg, accum_out_vec_2_msg, accum_out_vec_3_msg,
      accum_out_vec_4_msg, accum_out_vec_5_msg, accum_out_vec_6_msg, accum_out_vec_7_msg
);
  input clk;
  input rst;
  input write_req_val;
  output write_req_rdy;
  input [68:0] write_req_msg;
  input start_val;
  output start_rdy;
  input [5:0] start_msg;
  input weight_in_vec_0_val;
  input weight_in_vec_1_val;
  input weight_in_vec_2_val;
  input weight_in_vec_3_val;
  input weight_in_vec_4_val;
  input weight_in_vec_5_val;
  input weight_in_vec_6_val;
  input weight_in_vec_7_val;
  output weight_in_vec_0_rdy;
  output weight_in_vec_1_rdy;
  output weight_in_vec_2_rdy;
  output weight_in_vec_3_rdy;
  output weight_in_vec_4_rdy;
  output weight_in_vec_5_rdy;
  output weight_in_vec_6_rdy;
  output weight_in_vec_7_rdy;
  input [7:0] weight_in_vec_0_msg;
  input [7:0] weight_in_vec_1_msg;
  input [7:0] weight_in_vec_2_msg;
  input [7:0] weight_in_vec_3_msg;
  input [7:0] weight_in_vec_4_msg;
  input [7:0] weight_in_vec_5_msg;
  input [7:0] weight_in_vec_6_msg;
  input [7:0] weight_in_vec_7_msg;
  output accum_out_vec_0_val;
  output accum_out_vec_1_val;
  output accum_out_vec_2_val;
  output accum_out_vec_3_val;
  output accum_out_vec_4_val;
  output accum_out_vec_5_val;
  output accum_out_vec_6_val;
  output accum_out_vec_7_val;
  input accum_out_vec_0_rdy;
  input accum_out_vec_1_rdy;
  input accum_out_vec_2_rdy;
  input accum_out_vec_3_rdy;
  input accum_out_vec_4_rdy;
  input accum_out_vec_5_rdy;
  input accum_out_vec_6_rdy;
  input accum_out_vec_7_rdy;
  output [31:0] accum_out_vec_0_msg;
  output [31:0] accum_out_vec_1_msg;
  output [31:0] accum_out_vec_2_msg;
  output [31:0] accum_out_vec_3_msg;
  output [31:0] accum_out_vec_4_msg;
  output [31:0] accum_out_vec_5_msg;
  output [31:0] accum_out_vec_6_msg;
  output [31:0] accum_out_vec_7_msg;


  // Interconnect Declarations
  wire act_in_vec_0_val;
  wire act_in_vec_1_val;
  wire act_in_vec_2_val;
  wire act_in_vec_3_val;
  wire act_in_vec_4_val;
  wire act_in_vec_5_val;
  wire act_in_vec_6_val;
  wire act_in_vec_7_val;
  wire act_in_vec_0_rdy;
  wire act_in_vec_1_rdy;
  wire act_in_vec_2_rdy;
  wire act_in_vec_3_rdy;
  wire act_in_vec_4_rdy;
  wire act_in_vec_5_rdy;
  wire act_in_vec_6_rdy;
  wire act_in_vec_7_rdy;
  wire [7:0] act_in_vec_0_msg;
  wire [7:0] act_in_vec_1_msg;
  wire [7:0] act_in_vec_2_msg;
  wire [7:0] act_in_vec_3_msg;
  wire [7:0] act_in_vec_4_msg;
  wire [7:0] act_in_vec_5_msg;
  wire [7:0] act_in_vec_6_msg;
  wire [7:0] act_in_vec_7_msg;


  // Interconnect Declarations for Component Instantiations 
  SysArray sa_inst (
      .clk(clk),
      .rst(rst),
      .weight_in_vec_0_val(weight_in_vec_0_val),
      .weight_in_vec_1_val(weight_in_vec_1_val),
      .weight_in_vec_2_val(weight_in_vec_2_val),
      .weight_in_vec_3_val(weight_in_vec_3_val),
      .weight_in_vec_4_val(weight_in_vec_4_val),
      .weight_in_vec_5_val(weight_in_vec_5_val),
      .weight_in_vec_6_val(weight_in_vec_6_val),
      .weight_in_vec_7_val(weight_in_vec_7_val),
      .weight_in_vec_0_rdy(weight_in_vec_0_rdy),
      .weight_in_vec_1_rdy(weight_in_vec_1_rdy),
      .weight_in_vec_2_rdy(weight_in_vec_2_rdy),
      .weight_in_vec_3_rdy(weight_in_vec_3_rdy),
      .weight_in_vec_4_rdy(weight_in_vec_4_rdy),
      .weight_in_vec_5_rdy(weight_in_vec_5_rdy),
      .weight_in_vec_6_rdy(weight_in_vec_6_rdy),
      .weight_in_vec_7_rdy(weight_in_vec_7_rdy),
      .weight_in_vec_0_msg(weight_in_vec_0_msg),
      .weight_in_vec_1_msg(weight_in_vec_1_msg),
      .weight_in_vec_2_msg(weight_in_vec_2_msg),
      .weight_in_vec_3_msg(weight_in_vec_3_msg),
      .weight_in_vec_4_msg(weight_in_vec_4_msg),
      .weight_in_vec_5_msg(weight_in_vec_5_msg),
      .weight_in_vec_6_msg(weight_in_vec_6_msg),
      .weight_in_vec_7_msg(weight_in_vec_7_msg),
      .act_in_vec_0_val(act_in_vec_0_val),
      .act_in_vec_1_val(act_in_vec_1_val),
      .act_in_vec_2_val(act_in_vec_2_val),
      .act_in_vec_3_val(act_in_vec_3_val),
      .act_in_vec_4_val(act_in_vec_4_val),
      .act_in_vec_5_val(act_in_vec_5_val),
      .act_in_vec_6_val(act_in_vec_6_val),
      .act_in_vec_7_val(act_in_vec_7_val),
      .act_in_vec_0_rdy(act_in_vec_0_rdy),
      .act_in_vec_1_rdy(act_in_vec_1_rdy),
      .act_in_vec_2_rdy(act_in_vec_2_rdy),
      .act_in_vec_3_rdy(act_in_vec_3_rdy),
      .act_in_vec_4_rdy(act_in_vec_4_rdy),
      .act_in_vec_5_rdy(act_in_vec_5_rdy),
      .act_in_vec_6_rdy(act_in_vec_6_rdy),
      .act_in_vec_7_rdy(act_in_vec_7_rdy),
      .act_in_vec_0_msg(act_in_vec_0_msg),
      .act_in_vec_1_msg(act_in_vec_1_msg),
      .act_in_vec_2_msg(act_in_vec_2_msg),
      .act_in_vec_3_msg(act_in_vec_3_msg),
      .act_in_vec_4_msg(act_in_vec_4_msg),
      .act_in_vec_5_msg(act_in_vec_5_msg),
      .act_in_vec_6_msg(act_in_vec_6_msg),
      .act_in_vec_7_msg(act_in_vec_7_msg),
      .accum_out_vec_0_val(accum_out_vec_0_val),
      .accum_out_vec_1_val(accum_out_vec_1_val),
      .accum_out_vec_2_val(accum_out_vec_2_val),
      .accum_out_vec_3_val(accum_out_vec_3_val),
      .accum_out_vec_4_val(accum_out_vec_4_val),
      .accum_out_vec_5_val(accum_out_vec_5_val),
      .accum_out_vec_6_val(accum_out_vec_6_val),
      .accum_out_vec_7_val(accum_out_vec_7_val),
      .accum_out_vec_0_rdy(accum_out_vec_0_rdy),
      .accum_out_vec_1_rdy(accum_out_vec_1_rdy),
      .accum_out_vec_2_rdy(accum_out_vec_2_rdy),
      .accum_out_vec_3_rdy(accum_out_vec_3_rdy),
      .accum_out_vec_4_rdy(accum_out_vec_4_rdy),
      .accum_out_vec_5_rdy(accum_out_vec_5_rdy),
      .accum_out_vec_6_rdy(accum_out_vec_6_rdy),
      .accum_out_vec_7_rdy(accum_out_vec_7_rdy),
      .accum_out_vec_0_msg(accum_out_vec_0_msg),
      .accum_out_vec_1_msg(accum_out_vec_1_msg),
      .accum_out_vec_2_msg(accum_out_vec_2_msg),
      .accum_out_vec_3_msg(accum_out_vec_3_msg),
      .accum_out_vec_4_msg(accum_out_vec_4_msg),
      .accum_out_vec_5_msg(accum_out_vec_5_msg),
      .accum_out_vec_6_msg(accum_out_vec_6_msg),
      .accum_out_vec_7_msg(accum_out_vec_7_msg)
    );
  InputSetup is_inst (
      .clk(clk),
      .rst(rst),
      .write_req_val(write_req_val),
      .write_req_rdy(write_req_rdy),
      .write_req_msg(write_req_msg),
      .start_val(start_val),
      .start_rdy(start_rdy),
      .start_msg(start_msg),
      .act_in_vec_0_val(act_in_vec_0_val),
      .act_in_vec_1_val(act_in_vec_1_val),
      .act_in_vec_2_val(act_in_vec_2_val),
      .act_in_vec_3_val(act_in_vec_3_val),
      .act_in_vec_4_val(act_in_vec_4_val),
      .act_in_vec_5_val(act_in_vec_5_val),
      .act_in_vec_6_val(act_in_vec_6_val),
      .act_in_vec_7_val(act_in_vec_7_val),
      .act_in_vec_0_rdy(act_in_vec_0_rdy),
      .act_in_vec_1_rdy(act_in_vec_1_rdy),
      .act_in_vec_2_rdy(act_in_vec_2_rdy),
      .act_in_vec_3_rdy(act_in_vec_3_rdy),
      .act_in_vec_4_rdy(act_in_vec_4_rdy),
      .act_in_vec_5_rdy(act_in_vec_5_rdy),
      .act_in_vec_6_rdy(act_in_vec_6_rdy),
      .act_in_vec_7_rdy(act_in_vec_7_rdy),
      .act_in_vec_0_msg(act_in_vec_0_msg),
      .act_in_vec_1_msg(act_in_vec_1_msg),
      .act_in_vec_2_msg(act_in_vec_2_msg),
      .act_in_vec_3_msg(act_in_vec_3_msg),
      .act_in_vec_4_msg(act_in_vec_4_msg),
      .act_in_vec_5_msg(act_in_vec_5_msg),
      .act_in_vec_6_msg(act_in_vec_6_msg),
      .act_in_vec_7_msg(act_in_vec_7_msg)
    );
endmodule



